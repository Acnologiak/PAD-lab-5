��1     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.0.2�ub�n_estimators�K�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�auto�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Age��Sex��ChestPainType��	RestingBP��Cholesterol��	FastingBS��
RestingECG��MaxHR��ExerciseAngina��Oldpeak��ST_Slope�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h2�f8�����R�(KhONNNJ����J����K t�b�C              �?�t�bhSh&�scalar���hNC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hK�
node_count�KՌnodes�h(h+K ��h-��R�(KKՅ�h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hh2�i8�����R�(KhONNNJ����J����K t�bK ��h�h�K��h�h�K��h�h_K��h�h_K ��h�h�K(��h�h_K0��uK8KKt�b�B�.         T                    �?j8je3�?�           ��@                           �?���̟�?�            r@       
       
             �?X�If%��?\            �b@                           �?�Ru߬Α?G            �\@������������������������       �        4            �T@       	                    @K@      �?             @@                           f@P���Q�?             4@������������������������       �                     3@������������������������       �                     �?������������������������       �                     (@              	             �?�t����?             A@                           �?�z�G��?             $@                          �\@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                      @                           �?      �?             8@              	          ����?�}�+r��?
             3@                          �i@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@                           �L@���Q��?             @������������������������       �                      @������������������������       �                     @       C                    �?��t�?_            �a@       *                    @K@�e�}|�?N            �Z@       !       
             �? ����?0            @P@                           �I@@�E�x�?$            �H@������������������������       �                     E@                           `X@؇���X�?             @������������������������       �                     �?������������������������       �                     @"       )                    �?      �?             0@#       $                    �F@�q�q�?             "@������������������������       �                      @%       &                    �H@؇���X�?             @������������������������       �                     @'       (       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @+       @                    �?v�2t5�?            �D@,       3       
             �?^������?            �A@-       .                   Pc@���!pc�?             &@������������������������       �                     @/       2       	          ����?      �?             @0       1                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @4       ;                   �b@r�q��?             8@5       6                    `@P���Q�?             4@������������������������       �                     *@7       8       	          033�?؇���X�?             @������������������������       �                     @9       :                    �?      �?              @������������������������       �                     �?������������������������       �                     �?<       =                    �?      �?             @������������������������       �                      @>       ?                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?A       B                    _@r�q��?             @������������������������       �                     �?������������������������       �                     @D       O       	          @33�?">�֕�?            �A@E       J                    �?\X��t�?             7@F       G       
             �?X�Cc�?             ,@������������������������       �                     @H       I                   �`@      �?              @������������������������       �                     @������������������������       �                     @K       L                   �`@�����H�?             "@������������������������       �                     @M       N                   pa@      �?              @������������������������       �                     �?������������������������       �                     �?P       S                   �`@�8��8��?             (@Q       R                   �^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@U       �                    �?�����L�?           �{@V       �                    �?@�ܻ��?�            @u@W       �                   �f@^|�_��?\            �a@X                           �?
�K0��?Z             a@Y       n       
             �?�Gi����?G            �[@Z       i       	          ����?      �?!             H@[       b                     K@�ݜ�?            �C@\       a                   pf@�>����?             ;@]       `                   �[@ ��WV�?             :@^       _                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     7@������������������������       �                     �?c       h                   d@      �?	             (@d       e                    �?ףp=
�?             $@������������������������       �                     @f       g       	            �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @j       m                   `a@�<ݚ�?             "@k       l                   `U@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @o       |                    d@؇���X�?&            �O@p       q                    �K@�^����?#            �M@������������������������       �                     C@r       s                   �_@�q�q�?             5@������������������������       �                     @t       y                   0a@      �?             ,@u       v                   �`@؇���X�?             @������������������������       �                     @w       x       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?z       {       	          ����?؇���X�?             @������������������������       �                     �?������������������������       �                     @}       ~                   pn@      �?             @������������������������       �                      @������������������������       �                      @�       �       
             �?�	j*D�?             :@������������������������       �                     *@�       �                   �a@�n_Y�K�?             *@�       �       	             �?r�q��?             @������������������������       �                     @�       �                   Ps@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    @N@ ���3�?z            �h@�       �       
             �?X�If%��?Z            �b@�       �                   Pd@���Q��?
             .@�       �                    @M@      �?              @������������������������       �                     @�       �                    V@      �?             @�       �                   @X@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �b@���H��?P            �`@�       �                   `_@����y7�?L            @_@�       �                   �a@p��%���?,            @Q@�       �                    �?�:�^���?            �F@�       �                    a@Du9iH��?            �E@�       �                   0j@��?^�k�?            �A@�       �                   �X@�IєX�?
             1@������������������������       �                     �?������������������������       �        	             0@������������������������       �                     2@�       �                   �h@      �?              @������������������������       �                     @�       �                   �\@      �?             @������������������������       �                      @������������������������       �                      @�       �                     J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     8@�       �                   �\@؇���X�?              L@�       �                    �D@�q�q�?             5@������������������������       �                     @�       �                   �m@��S���?             .@�       �                   0i@�<ݚ�?             "@������������������������       �                     @�       �                   �b@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �       	          ����?��?^�k�?            �A@�       �                   �`@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     <@�       �                    q@      �?              @�       �                   c@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    �?p���?              I@������������������������       �                     >@�       �                   �a@P���Q�?             4@������������������������       �                     0@�       �                   p@      �?             @������������������������       �                     �?������������������������       �                     @�       �       
             �? >�֕�?@            @Z@�       �                   `\@      �?	             (@������������������������       �                     @�       �                   @b@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   ``@�g�y��?7            @W@������������������������       �                     E@�       �                   �`@�IєX�?            �I@������������������������       �                      @�       �       	          `ff�?@�E�x�?            �H@������������������������       �                     B@�       �                   @^@$�q-�?             *@�       �                    �?r�q��?             @�       �                    �Q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�b�values�h(h+K ��h-��R�(KK�KK��h_�BP       Ps@     �z@      j@      T@     �^@      9@     @\@      �?     �T@              ?@      �?      3@      �?      3@                      �?      (@              $@      8@      @      @      @      �?              �?      @                       @      @      5@      �?      2@      �?      @      �?                      @              (@       @      @       @                      @     �U@     �K@     �R@      ?@      M@      @      H@      �?      E@              @      �?              �?      @              $@      @      @      @       @              �?      @              @      �?      �?              �?      �?              @              1@      8@      (@      7@       @      @      @              �?      @      �?      �?      �?                      �?               @      @      4@      �?      3@              *@      �?      @              @      �?      �?      �?                      �?      @      �?       @              �?      �?      �?                      �?      @      �?              �?      @              &@      8@      $@      *@      "@      @      @              @      @      @                      @      �?       @              @      �?      �?      �?                      �?      �?      &@      �?      �?              �?      �?                      $@      Y@     �u@     �W@     �n@      Q@     �R@     �O@     �R@     �F@     �P@      B@      (@      A@      @      9@       @      9@      �?       @      �?       @                      �?      7@                      �?      "@      @      "@      �?      @              @      �?      @                      �?               @       @      @       @      �?              �?       @                      @      "@      K@      @      J@              C@      @      ,@              @      @      @      @      �?      @               @      �?       @                      �?      �?      @      �?                      @       @       @       @                       @      2@       @      *@              @       @      @      �?      @               @      �?       @                      �?              @      @              :@     �e@      9@     �^@      "@      @       @      @              @       @       @       @      �?              �?       @                      �?      @              0@     @]@      (@     @\@      @     @P@      @     �D@      @      D@      �?      A@      �?      0@      �?                      0@              2@       @      @              @       @       @       @                       @      �?      �?      �?                      �?              8@       @      H@      @      ,@              @      @       @      @       @      @              @       @      @                       @              @      �?      A@      �?      @      �?                      @              <@      @      @       @      @       @                      @       @              �?     �H@              >@      �?      3@              0@      �?      @      �?                      @      @     �X@      @      "@              @      @       @      @                       @      @     �V@              E@      @      H@       @              �?      H@              B@      �?      (@      �?      @      �?      �?              �?      �?                      @              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKᅔh~�B81         X       
             �?4�5����?�           ��@       #                    �?`}�?��?�            �t@                          �P@���ۑ��?x            �h@                           �?և���X�?             ,@                           �?���!pc�?             &@������������������������       �                      @������������������������       �                     @������������������������       �                     @	                           @L@@-�_ .�?p             g@
                          �g@pY���D�?`            �c@                          @[@ u�z\A�?_            `c@                           @G@�C��2(�?             &@������������������������       �                      @                           �?�q�q�?             @������������������������       �                     �?                          `m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        Y             b@������������������������       �                     @       "                    �?�<ݚ�?             ;@                          Pc@���Q��?
             .@                           �?z�G�z�?             $@                          �`@�q�q�?             @                          @b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @       !                    �N@z�G�z�?             @               	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     (@$       O                    �?�c��{-�?P            ``@%       >                    �?���I���?A            �[@&       9       	          ����?ޭ�W[��?,            @T@'       4                    �L@��ɉ�?"            @P@(       /                    ]@���}<S�?             G@)       .                   �p@      �?             (@*       -                   i@ףp=
�?             $@+       ,                   �X@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @0       1                   �b@г�wY;�?             A@������������������������       �                     @@2       3                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?5       8                   �b@�d�����?	             3@6       7                   @q@@�0�!��?             1@������������������������       �                     ,@������������������������       �                     @������������������������       �                      @:       ;                    �J@      �?
             0@������������������������       �                     @<       =                    a@���Q��?             $@������������������������       �                     @������������������������       �                     @?       N                    c@d��0u��?             >@@       M                    �?R�}e�.�?             :@A       L       	          033�?�+e�X�?             9@B       G                    �I@�����?             3@C       F                   �`@����X�?             @D       E       	          `ff�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @H       K                    �N@�8��8��?             (@I       J                   �b@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @P       U                   ``@R���Q�?             4@Q       R                    ]@      �?             0@������������������������       �        	             ,@S       T                   �]@      �?              @������������������������       �                     �?������������������������       �                     �?V       W       	          433�?      �?             @������������������������       �                      @������������������������       �                      @Y       �                    �?P� �&�?           @y@Z       �                    �?BgG�".�?�            `q@[       �                   P`@8�ƨxt�?�            �k@\       m                    �?     8�?S             `@]       d                    @H@ҳ�wY;�?             A@^       _                   �[@X�Cc�?	             ,@������������������������       �                     @`       c                   Pd@"pc�
�?             &@a       b                   �c@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @e       j                   �d@R���Q�?             4@f       g                   �m@�����H�?             2@������������������������       �                     .@h       i                   �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @k       l                    �?      �?              @������������������������       �                     �?������������������������       �                     �?n       �                   0a@�*/�8V�?:            �W@o       v                    @L@����p�?+             Q@p       q                    �? ���J��?            �C@������������������������       �                     9@r       u                   �\@@4և���?
             ,@s       t       	              @z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@w       z                    �L@\-��p�?             =@x       y                   �d@�q�q�?             @������������������������       �                     �?������������������������       �                      @{       �                    �?$�q-�?             :@|                           @P@r�q��?             @}       ~                     O@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       	          ����?P���Q�?             4@������������������������       �                     �?������������������������       �        
             3@�       �                    �?���B���?             :@�       �       	             �?�IєX�?
             1@������������������������       �                     &@�       �       	             @r�q��?             @�       �                   @Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    ^@X�<ݚ�?             "@�       �                   �a@z�G�z�?             @�       �                   �n@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �? rpa�?B            @W@�       �                    �?      �?             0@�       �                    �?      �?              @������������������������       �                     �?�       �                    �K@؇���X�?             @������������������������       �                     @�       �                    a@�q�q�?             @������������������������       �                     �?�       �                   �i@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   n@      �?              @������������������������       �                      @������������������������       �                     @�       �                   �a@�e���@�?6            @S@�       �       	             �?г�wY;�?             A@�       �       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     ?@������������������������       �                    �E@�       �                   a@�^���U�?$            �L@�       �                   �Q@\-��p�?             =@������������������������       �                     �?�       �                    Z@ �Cc}�?             <@������������������������       �                      @�       �                    �? ��WV�?             :@������������������������       �        
             1@�       �                    @K@�����H�?             "@�       �                   0a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?X�Cc�?             <@�       �                   @\@և���X�?             @������������������������       �                     �?�       �                   Pc@�q�q�?             @������������������������       �                     @�       �       	          033�?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	          ����?����X�?             5@�       �                   0c@X�<ݚ�?             "@�       �       	          433�?�q�q�?             @������������������������       �                     �?�       �                   @b@���Q��?             @������������������������       �                      @�       �                    �H@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?�8��8��?             (@�       �       	          `ff@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �c@�����?H            �_@�       �                   pb@ '��h�?A            @[@�       �                   �Q@�}��L�?+            �R@�       �                   �l@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        )            @R@�       �                   P`@�t����?             A@�       �                   �[@���7�?             6@������������������������       �                     &@�       �                    ]@�C��2(�?             &@�       �                   @p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                   Pa@      �?             (@�       �                   �j@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   @d@j���� �?             1@������������������������       �                     @������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KK�KK��h_�B       �t@     y@     0p@     �Q@     �f@      0@       @      @       @      @       @                      @              @     �e@      $@     @c@      @     @c@      �?      $@      �?       @               @      �?      �?              �?      �?      �?                      �?      b@                      @      5@      @      "@      @       @       @      @       @      �?       @               @      �?              @              @              �?      @      �?       @      �?                       @               @      (@              S@     �K@     @R@      C@      O@      3@      L@      "@      E@      @      "@      @      "@      �?      �?      �?      �?                      �?       @                       @     �@@      �?      @@              �?      �?      �?                      �?      ,@      @      ,@      @      ,@                      @               @      @      $@              @      @      @              @      @              &@      3@      @      3@      @      3@      @      *@      @       @      �?       @               @      �?              @              �?      &@      �?      @              @      �?                       @              @      �?              @              @      1@      �?      .@              ,@      �?      �?      �?                      �?       @       @       @                       @     �R@     �t@      O@      k@      ;@     @h@      6@     �Z@      (@      6@      "@      @              @      "@       @       @       @       @                       @      @              @      1@       @      0@              .@       @      �?              �?       @              �?      �?      �?                      �?      $@      U@      @     �O@      �?      C@              9@      �?      *@      �?      @              @      �?                      "@      @      9@       @      �?              �?       @               @      8@      �?      @      �?      �?              �?      �?                      @      �?      3@      �?                      3@      @      5@      �?      0@              &@      �?      @      �?       @      �?                       @              @      @      @      @      �?       @      �?       @                      �?       @                      @      @      V@      @      (@       @      @      �?              �?      @              @      �?       @              �?      �?      �?      �?                      �?       @      @       @                      @      �?      S@      �?     �@@      �?       @               @      �?                      ?@             �E@     �A@      6@      9@      @              �?      9@      @               @      9@      �?      1@               @      �?       @      �?              �?       @              @              $@      2@      @      @              �?      @       @      @              �?       @               @      �?              @      .@      @      @       @      @              �?       @      @               @       @      �?       @                      �?      @              �?      &@      �?      @              @      �?                      @      (@     �\@      @      Z@      �?     �R@      �?      �?              �?      �?                     @R@      @      >@      �?      5@              &@      �?      $@      �?      �?              �?      �?                      "@      @      "@      @       @               @      @                      @      @      $@      @                      $@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKׅ�h~�B/         ^       	          ����?p�Vv���?�           ��@       ?                    �?X~�pX��?�            �v@       &       
             �?BA�V�?�            �r@                          �b@ d�=��?�            @l@                          �O@X�?٥�?�            �i@                           �?�eP*L��?             &@������������������������       �                     @������������������������       �                     @	              	            �? ���J��?z            `h@
                          Pb@ }�Я��?p            @f@                          �[@ A��� �?g            @d@                          �h@ �q�q�?             8@                            G@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     3@������������������������       �        Y            @a@                          �d@      �?	             0@                          �b@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@                          �a@@�0�!��?
             1@������������������������       �                     "@                          �a@      �?              @������������������������       �                      @              	            �?r�q��?             @������������������������       �                     @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?        #                   �c@�z�G��?             4@!       "                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @$       %                   �g@@4և���?	             ,@������������������������       �                     *@������������������������       �                     �?'       (                   �`@      �?0             R@������������������������       �                     1@)       2                    �?��N`.�?#            �K@*       +                    �D@V������?            �B@������������������������       �                     $@,       1                    �?�5��?             ;@-       0                   pm@z�G�z�?             4@.       /       	          ����?���Q��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     $@������������������������       �                     @3       >                   �q@b�2�tk�?             2@4       7                   @k@      �?             ,@5       6                   �h@z�G�z�?             @������������������������       �                     �?������������������������       �                     @8       =                   @a@�q�q�?             "@9       <                    �?���Q��?             @:       ;                   �c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @@       E                    ]@��y�:�?,            �P@A       D                    �?      �?              @B       C                    �D@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @F       ]                   Pd@�k��(A�?&            �M@G       X                    �?���B���?"             J@H       U                   �s@�˹�m��?             C@I       P       	          ����?�X�<ݺ?             B@J       K                   pb@(;L]n�?             >@������������������������       �                     9@L       O                     K@z�G�z�?             @M       N                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @Q       T                    [@r�q��?             @R       S                   p`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @V       W                   �t@      �?              @������������������������       �                     �?������������������������       �                     �?Y       Z                    �?      �?             ,@������������������������       �                     @[       \                   �b@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @_       ~       
             �?�zц��?�            w@`       u                    �?�g�y��?(             O@a       b                   �^@4�B��?            �B@������������������������       �                     @c       t                   `f@     ��?             @@d       m                    �L@r�q��?             >@e       f                    �?�}�+r��?             3@������������������������       �                     &@g       l                   �j@      �?              @h       k                    �?�q�q�?             @i       j                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @n       o                    a@���|���?             &@������������������������       �                     @p       q       	          ����?      �?              @������������������������       �                     @r       s                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @v       w                   �Y@z�G�z�?             9@������������������������       �                     @x       }       	          `ff�?���N8�?             5@y       z                    �?z�G�z�?             @������������������������       �                     @{       |                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             0@       �                    �?/ĕn�?�            0s@�       �                   �s@lutee�?.            �P@�       �                   �c@     x�?,             P@�       �                    �?�*/�8V�?!            �G@�       �       	          `ff�?     ��?             @@�       �                   �[@��S���?             .@������������������������       �                     @�       �                   @c@�q�q�?
             (@�       �                    ^@z�G�z�?             $@������������������������       �                     @�       �                   �`@����X�?             @������������������������       �                     �?�       �                   @_@r�q��?             @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                   m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    b@�t����?	             1@�       �                   @a@���Q��?             @������������������������       �                      @�       �                   Pn@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@�       �                    �?�r����?             .@�       �       	             �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     $@�       �                   �\@ҳ�wY;�?             1@������������������������       �                     @�       �                   pe@d}h���?	             ,@�       �                   (p@8�Z$���?             *@������������������������       �                     &@������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �Q@��(\���?�             n@�       �                   pb@�j�-��?�            `l@�       �       	          ����?�F�l���?�            �g@�       �                    �L@,���i�?            �D@�       �                    @L@�E��ӭ�?             2@�       �                    �?     ��?             0@�       �                   �l@@4և���?             ,@������������������������       �                     $@�       �                   p@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     7@�       �                   �_@p���?i            �b@�       �       	          033�?Du9iH��?            �E@������������������������       �                     *@�       �                    �?ףp=
�?             >@�       �                   @M@�����H�?             ;@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       	          ����?�8��8��?             8@�       �                    �G@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    p@���7�?             6@������������������������       �                     ,@�       �                    �J@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        J            �Z@�       �                   �a@r�q��?             B@�       �       	          033�?V�a�� �?             =@�       �                    �N@�}�+r��?             3@������������������������       �                     ,@�       �                    @O@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    @N@      �?             $@�       �                   �d@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   `@�	j*D�?             *@������������������������       �                     @������������������������       �                     "@�t�bh�h(h+K ��h-��R�(KK�KK��h_�Bp       @t@     �y@     @o@     �\@     �l@     �Q@     @j@      0@     �h@      $@      @      @      @                      @     �g@      @      f@       @      d@      �?      7@      �?      @      �?              �?      @              3@             @a@              .@      �?      @      �?              �?      @              "@              ,@      @      "@              @      @               @      @      �?      @              �?      �?      �?                      �?      ,@      @      �?      @      �?                      @      *@      �?      *@                      �?      2@      K@              1@      2@     �B@      &@      :@              $@      &@      0@      @      0@      @      @              @      @                      $@      @              @      &@      @      @      �?      @      �?                      @      @      @       @      @       @      �?       @                      �?               @      @                      @      6@     �F@      @      @       @      @       @                      @      @              1@      E@      $@      E@      @     �A@       @      A@      �?      =@              9@      �?      @      �?      �?              �?      �?                      @      �?      @      �?       @               @      �?                      @      �?      �?      �?                      �?      @      @      @               @      @              @       @              @             �R@     pr@      >@      @@      9@      (@              @      9@      @      9@      @      2@      �?      &@              @      �?       @      �?      �?      �?              �?      �?              �?              @              @      @              @      @      �?      @               @      �?       @                      �?               @      @      4@      @              �?      4@      �?      @              @      �?      �?              �?      �?                      0@      F@     pp@      :@     �D@      7@     �D@      (@     �A@      $@      6@       @      @              @       @      @       @       @      @              @       @              �?      @      �?       @      �?      �?              �?      �?      �?                      �?      @                       @       @      .@       @      @               @       @      �?       @                      �?              (@       @      *@       @      @       @                      @              $@      &@      @              @      &@      @      &@       @      &@                       @              �?      @              2@     �k@      ,@     �j@       @     �f@      @      B@      @      *@      @      *@      �?      *@              $@      �?      @      �?                      @       @               @                      7@      @     `b@      @      D@              *@      @      ;@      @      8@      �?       @      �?                       @       @      6@      �?      �?              �?      �?              �?      5@              ,@      �?      @      �?                      @              @             �Z@      @      >@      @      7@      �?      2@              ,@      �?      @      �?                      @      @      @      @       @      @                       @              @              @      @      "@      @                      "@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKׅ�h~�B/         t                    �?U�ք�?�           ��@       3                    �?n�����?           @z@              
             �?�R�� �?�             n@                          �O@H��2�?z            @g@                           �N@X�<ݚ�?             "@������������������������       �                     @                           ^@r�q��?             @������������������������       �                     @	       
                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                          h@���fG��?s             f@                           �O@�C��2(�?r             f@              	          ���@ t�)Ї?o            `e@������������������������       �        n            @e@������������������������       �                     �?                          @t@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?                           �a@�eP*L��?(            �K@                          �`@z�G�z�?             4@                           �?���|���?             &@                           �?؇���X�?             @                          @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                          �m@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@!       .                    �?���Q��?            �A@"       #                     G@�ՙ/�?             5@������������������������       �                     @$       -                    �?�E��ӭ�?             2@%       ,                    �?     ��?             0@&       +                   �p@���Q��?             @'       *                   Pm@      �?             @(       )       	          hff�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     &@������������������������       �                      @/       2                    �H@@4և���?
             ,@0       1                   d@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@4       =                   @E@���i!��?u            `f@5       <                    �?@4և���?             E@6       ;                   �^@      �?             @7       :                   `]@      �?             @8       9                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     B@>       Y                    �J@���<��?Y             a@?       B                    a@H(���o�?%            �J@@       A       
             �?�q�q�?
             (@������������������������       �                     @������������������������       �                     @C       F                    @D@������?            �D@D       E                    �?      �?              @������������������������       �                     @������������������������       �                      @G       R       
             �?"pc�
�?            �@@H       Q       	          ����?$�q-�?             :@I       J                    �?�C��2(�?             6@������������������������       �        	             ,@K       L                   0j@      �?              @������������������������       �                     �?M       N                   Pb@؇���X�?             @������������������������       �                     @O       P                    p@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @S       T                   `]@և���X�?             @������������������������       �                     �?U       V       	          ����?�q�q�?             @������������������������       �                     @W       X                    @I@�q�q�?             @������������������������       �                     �?������������������������       �                      @Z       e       
             �?�q�q�?4             U@[       `                   Po@���N8�?             5@\       ]                    b@��S�ۿ?             .@������������������������       �        
             *@^       _       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?a       d                    @M@�q�q�?             @b       c                   �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @f       i       	          ����?��s����?#            �O@g       h       	          833�?�LQ�1	�?             7@������������������������       �                     .@������������������������       �                      @j       o                    `P@ףp=
�?             D@k       n                    @M@ >�֕�?            �A@l       m       	             �?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @������������������������       �                     :@p       s                    �?���Q��?             @q       r                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @u       �       
             �?JN�#:�?�            �s@v       {                    I@\X��t�?             G@w       x                   b@�C��2(�?             &@������������������������       �                     "@y       z                    �K@      �?              @������������������������       �                     �?������������������������       �                     �?|       �                    `@����X�?            �A@}       �       	          ����?��
ц��?             *@~                           �?      �?              @������������������������       �                     @������������������������       �                     @�       �                   �a@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �       	          033�?"pc�
�?             6@������������������������       �                     0@�       �                    �H@�q�q�?             @������������������������       �                      @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �                   P`@pH����?�            �p@�       �       	          ����?b�h�d.�?I            @Z@�       �                   0a@j�g�y�?-             O@�       �                    @L@(L���?"            �E@�       �                   ps@���7�?             6@������������������������       �                     2@�       �                   �t@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �d@���N8�?             5@������������������������       �        	             (@�       �                   xt@X�<ݚ�?             "@�       �                    �N@����X�?             @������������������������       �                     @�       �                   (p@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    �?�\��N��?             3@�       �                    �?"pc�
�?             &@�       �       	             �?      �?              @�       �                   `h@�q�q�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   �Z@Du9iH��?            �E@�       �                   �X@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?P���Q�?             D@������������������������       �                     6@�       �                   �a@�����H�?             2@�       �                   @\@�IєX�?             1@�       �                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        
             ,@������������������������       �                     �?�       �                    �?��|r�{�?b            `d@�       �                   @s@PX�V|�?S            `a@�       �                   `f@�i�y�?K            �_@�       �       	          ����? ����?F            �]@�       �                   �`@�7��?            �C@�       �                    �?�?�|�?            �B@������������������������       �                      @�       �                    �K@��?^�k�?            �A@�       �                   �\@      �?              @�       �                    �I@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     ;@�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        0             T@�       �                    �?����X�?             @������������������������       �                     �?�       �                    �?�q�q�?             @�       �                    a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?�θ�?             *@������������������������       �                     "@�       �       	             �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �a@      �?             8@������������������������       �                     "@�       �                    �?z�G�z�?	             .@������������������������       �                     @������������������������       �                     (@�t�bh�h(h+K ��h-��R�(KK�KK��h_�Bp        t@     �y@     �p@      c@     `i@      C@     @f@       @      @      @              @      @      �?      @               @      �?       @                      �?     �e@      @     �e@      @     @e@      �?     @e@                      �?      @       @      @                       @              �?      9@      >@      @      0@      @      @      �?      @      �?      �?              �?      �?                      @      @      �?      @                      �?              "@      5@      ,@       @      *@      @              @      *@      @      *@      @       @      @      �?      �?      �?      �?                      �?       @                      �?              &@       @              *@      �?      @      �?              �?      @              "@             @P@     �\@      @     �C@      @      @      @      �?      �?      �?      �?                      �?       @                       @              B@      O@     �R@      A@      3@      @      @      @                      @      =@      (@       @      @              @       @              ;@      @      8@       @      4@       @      ,@              @       @              �?      @      �?      @               @      �?       @                      �?      @              @      @      �?               @      @              @       @      �?              �?       @              <@      L@      0@      @      ,@      �?      *@              �?      �?              �?      �?               @      @       @      �?       @                      �?              @      (@     �I@       @      .@              .@       @              @      B@       @     �@@       @      @       @                      @              :@       @      @       @      �?              �?       @                       @      K@     @p@      :@      4@      �?      $@              "@      �?      �?              �?      �?              9@      $@      @      @      @      @      @                      @      @      �?      @                      �?      2@      @      0@               @      @               @       @       @               @       @              <@      n@      2@     �U@      .@     �G@      @     �B@      �?      5@              2@      �?      @      �?                      @      @      0@              (@      @      @      @       @      @              �?       @               @      �?                       @      "@      $@      "@       @      @       @      �?       @              �?      �?      �?      �?                      �?      @              @                       @      @      D@      �?       @               @      �?               @      C@              6@       @      0@      �?      0@      �?       @               @      �?                      ,@      �?              $@      c@      @     �`@      @     �^@       @     @]@       @     �B@      �?      B@               @      �?      A@      �?      @      �?       @               @      �?                      @              ;@      �?      �?      �?                      �?              T@       @      @              �?       @      @       @      �?       @                      �?              @      @      $@              "@      @      �?              �?      @              @      5@              "@      @      (@      @                      (@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKㅔh~�B�1         L                    �?4�5����?�           ��@       A                    �?Z�/�j��?�            �r@       (                    @L@T$�#���?�            `n@              
             �?��H���?|             h@                          �g@P�Lt�<�?d             c@                          pf@�}��L�?c            �b@                           �?���б�?X            �`@       	                   @n@�����?D            @Y@������������������������       �        (             M@
                          0c@ qP��B�?            �E@                          �n@      �?
             0@������������������������       �                     �?������������������������       �        	             .@������������������������       �                     ;@������������������������       �                     A@                           �?��S�ۿ?             .@������������������������       �                     &@                          �`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @       '                   0a@��]�T��?            �D@       &                    �?�E��ӭ�?             B@       %                    �?�eP*L��?             6@                            �?�\��N��?             3@                           @C@���|���?             &@������������������������       �                     @              	          033�?�q�q�?             @������������������������       �                     @                          �i@�q�q�?             @������������������������       �                     �?������������������������       �                      @!       $                    �?      �?              @"       #                   �r@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     ,@������������������������       �                     @)       ,                    �?��H�}�?$             I@*       +                    _@8�Z$���?
             *@������������������������       �                      @������������������������       �        	             &@-       .                   `\@��J�fj�?            �B@������������������������       �                     @/       0                   �^@���|���?            �@@������������������������       �                      @1       <       	          ����?�q�����?             9@2       3                   �`@p�ݯ��?             3@������������������������       �                      @4       ;       	          ����?�t����?             1@5       :                   �d@�eP*L��?             &@6       7                   �j@      �?              @������������������������       �                     @8       9                   `c@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @=       >                    �?r�q��?             @������������������������       �                     @?       @                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?B       C                    �G@��N`.�?'            �K@������������������������       �                     @D       E                   �]@ \� ���?#            �H@������������������������       �                     1@F       G       
             �?      �?             @@������������������������       �                     "@H       K                    �?�LQ�1	�?             7@I       J                   �s@���N8�?             5@������������������������       �                     4@������������������������       �                     �?������������������������       �                      @M       �       	          ����?      �?           @{@N       w       
             �?\`*�s�?k             e@O       p                    �?�
�G�?6             V@P       ]                    �?�sly47�?/            �R@Q       R                   @^@      �?             @@������������������������       �        	             *@S       \                    �?���y4F�?             3@T       [                    @N@�	j*D�?	             *@U       V                    W@      �?             (@������������������������       �                      @W       X                   `k@ףp=
�?             $@������������������������       �                     @Y       Z                   @b@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @^       m                    b@�+��<��?            �E@_       l                   pf@��.k���?             A@`       e                   �`@X�Cc�?             <@a       d                   @Y@�q�q�?             (@b       c                   �[@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @f       g                    @H@      �?	             0@������������������������       �                     $@h       k                    �?�q�q�?             @i       j                    �N@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @n       o                   pc@�����H�?             "@������������������������       �                      @������������������������       �                     �?q       v                   ``@��
ц��?             *@r       u                     K@�q�q�?             "@s       t                   �[@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @x       y                   �g@z�G�z�?5             T@������������������������       �                     B@z       {                   �_@�X����?             F@������������������������       �                     0@|       �                     P@      �?             <@}       �                   �p@�ՙ/�?             5@~       �                    �?�E��ӭ�?             2@       �                   �m@�eP*L��?	             &@�       �                    `@����X�?             @������������������������       �                     �?�       �                   @l@r�q��?             @�       �                    @N@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       	          ����?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                   �`@��v����?�            �p@�       �                    �?V�a�� �?L             ]@�       �                   �j@ܩ�d	��?4            �S@�       �                    Y@��
ц��?             :@������������������������       �                     @�       �                    @I@�û��|�?             7@�       �                   �Z@ףp=
�?             $@�       �                    �D@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   `i@�n_Y�K�?	             *@�       �       	             �?���!pc�?             &@������������������������       �                      @�       �                    �?�����H�?             "@������������������������       �                     @�       �                   �f@z�G�z�?             @������������������������       �                     @�       �                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �e@�iʫ{�?#            �J@�       �       	          ����?8��8���?!             H@�       �                    �?z�G�z�?             4@�       �                    �H@      �?
             0@�       �                    �F@���Q��?             @������������������������       �                      @�       �                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@�       �                   �`@      �?             @������������������������       �                      @������������������������       �                      @�       �       	          ���@h�����?             <@������������������������       �                     7@�       �                   �r@z�G�z�?             @�       �                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   `]@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   �x@�L���?            �B@�       �       
             �?��?^�k�?            �A@�       �       	          033�?�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     :@������������������������       �                      @�       �                    �R@�˹�m��?e             c@�       �                   �b@@�+9\J�?d            �b@�       �                    `P@Pa�	�?S            �`@�       �       	          ����?0�)AU��?J            �\@�       �                    �? �q�q�?!             H@������������������������       �                     ;@�       �                   �_@�����?             5@������������������������       �                     0@�       �       
             �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �        )            �P@�       �       	          033@�����H�?	             2@������������������������       �                     $@�       �                     Q@      �?              @������������������������       �                      @������������������������       �                     @�       �                    �?p�ݯ��?             3@�       �       	          `ff@��
ц��?             *@�       �                    �F@�q�q�?	             "@������������������������       �                      @�       �       	          033�?և���X�?             @�       �                   �d@���Q��?             @�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �       
             �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�t�b��     h�h(h+K ��h-��R�(KK�KK��h_�B0       �t@     y@      l@     �R@     �i@     �B@     �e@      3@     �b@      @     �b@       @     �`@      �?      Y@      �?      M@              E@      �?      .@      �?              �?      .@              ;@              A@              ,@      �?      &@              @      �?              �?      @                       @      :@      .@      :@      $@      (@      $@      "@      $@      @      @              @      @       @      @              �?       @      �?                       @      @      @      �?      @              @      �?              @              @              ,@                      @      @@      2@      &@       @               @      &@              5@      0@              @      5@      (@       @              *@      (@      (@      @               @      (@      @      @      @      @      @              @      @       @      @                       @      @              @              �?      @              @      �?       @               @      �?              2@     �B@      @              (@     �B@              1@      (@      4@      "@              @      4@      �?      4@              4@      �?               @             @[@     pt@     @R@     �W@     �M@      =@      J@      7@      <@      @      *@              .@      @      "@      @      "@      @               @      "@      �?      @              @      �?      @                      �?              �?      @              8@      3@      0@      2@      $@      2@       @      @       @      @              @       @              @               @      ,@              $@       @      @       @       @       @                       @               @      @               @      �?       @                      �?      @      @      @      @      @       @      @                       @              @      @              ,@     �P@              B@      ,@      >@              0@      ,@      ,@      *@       @      *@      @      @      @      @       @              �?      @      �?       @      �?       @                      �?      @              �?      @      �?                      @      @                      @      �?      @              @      �?              B@      m@      8@      W@      5@      M@      (@      ,@      @              "@      ,@      �?      "@      �?      �?              �?      �?                       @       @      @       @      @               @       @      �?      @              @      �?      @              �?      �?              �?      �?                       @      "@      F@      @     �E@      @      0@       @      ,@       @      @               @       @      �?              �?       @                      &@       @       @       @                       @      �?      ;@              7@      �?      @      �?       @      �?                       @               @      @      �?      @                      �?      @      A@      �?      A@      �?       @      �?                       @              :@       @              (@     �a@      &@     �a@      @      `@       @      \@       @      G@              ;@       @      3@              0@       @      @       @                      @             �P@       @      0@              $@       @      @       @                      @      @      (@      @      @      @      @       @              @      @       @      @       @      �?       @                      �?               @       @                      @      �?      @      �?                      @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B8*         V       	          ����?6������?�           ��@       =       
             �?��_���?�             w@                          @E@(��R%��?�            �p@                          �[@��H�}�?             9@������������������������       �                     @                           �?�\��N��?             3@                           �?���Q��?	             .@                           �?      �?             (@	       
       	          hff�?�����H�?             "@������������������������       �                      @������������������������       �                     �?                          �]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @       <                    �R@�l�T{�?�             n@                          �b@x�U���?�            �m@                          Hp@ ����?L            �]@������������������������       �        :             X@                          �b@���}<S�?             7@                           _@���N8�?             5@                          �^@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     0@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?       #                   0c@�r����?O             ^@       "                    �?z�G�z�?             @        !                   c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @$       7                    b@������?L            �\@%       ,                    �L@����?E            @Z@&       '                    �?����?�?;            �V@������������������������       �        0             S@(       +                     E@؇���X�?             ,@)       *                   `d@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     "@-       6                    �?���Q��?
             .@.       5                    �?���Q��?             $@/       0                   �`@      �?              @������������������������       �                     @1       2                   @f@      �?             @������������������������       �                     �?3       4                   `q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @8       ;                   �c@���Q��?             $@9       :                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @>       ?                   ph@�4�M�f�?@            �Y@������������������������       �                     D@@       C                    �?V��z4�?%             O@A       B                    �?���|���?             &@������������������������       �                     @������������������������       �                     @D       S                    �O@������?            �I@E       H                   �h@      �?             D@F       G       	          ����?���Q��?             @������������������������       �                      @������������������������       �                     @I       N       	          ����? >�֕�?            �A@J       K                   pe@      �?             @@������������������������       �                     ;@L       M                    �F@z�G�z�?             @������������������������       �                     �?������������������������       �                     @O       R                    �?�q�q�?             @P       Q                    �K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?T       U       	          ����?���|���?             &@������������������������       �                     @������������������������       �                     @W       �                   �`@xƅd�?�            �v@X       y       	          pff�?ܷ��?��?~            `i@Y       r                    �?4Ky\�?L            @\@Z       e                    �?8EGr��?B             Y@[       d       	          ����?�q�q�?             8@\       _                    �?�GN�z�?             6@]       ^                   �v@      �?              @������������������������       �                     @������������������������       �                      @`       c                   �`@d}h���?	             ,@a       b                   �^@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@������������������������       �                      @f       q                    �?�}�+r��?2             S@g       h                    _@ 	��p�?%             M@������������������������       �                    �E@i       j       
             �?������?             .@������������������������       �                      @k       l                     L@8�Z$���?	             *@������������������������       �                     "@m       n                   @Z@      �?             @������������������������       �                     �?o       p                    �M@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     2@s       t       	          pff�?��
ц��?
             *@������������������������       �                     @u       x                   �f@      �?              @v       w                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @z       {       	          `ff@`Ӹ����?2            �V@������������������������       �        $            �P@|       �                    �?r�q��?             8@}       �                    �J@��2(&�?             6@~                          �`@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �        	             1@�       �                   Hq@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ���@噼:��?d            `d@�       �                   `U@:��au��?I            �^@�       �       	          ����?�<ݚ�?             2@������������������������       �                     (@�       �                   �b@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �M@&RN���?>            @Z@�       �                    �?      �?/             T@�       �                   �[@���H��?             E@������������������������       �                      @�       �                    �L@��(\���?             D@������������������������       �                    �A@�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   0c@P����?             C@�       �                   �a@R���Q�?             4@�       �                    �J@      �?              @�       �                    �E@r�q��?             @������������������������       �                     @�       �                    a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     (@�       �                   q@X�<ݚ�?
             2@�       �                   0i@�z�G��?             $@������������������������       �                     @������������������������       �                     @�       �                    �?      �?              @�       �                   �q@z�G�z�?             @������������������������       �                      @�       �                   �r@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �n@`�Q��?             9@�       �                    e@      �?              @�       �                    �P@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �       	          ����?@�0�!��?	             1@������������������������       �                     @������������������������       �                     ,@�       �                   �j@��(\���?             D@�       �                    Z@8�Z$���?	             *@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@�       �                   ``@ 7���B�?             ;@�       �                    �?�����H�?             "@�       �                    n@r�q��?             @������������������������       �                     @�       �                   �e@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     2@�t�bh�h(h+K ��h-��R�(KK�KK��h_�B       �t@     �x@      o@     �]@     �l@      B@      "@      0@              @      "@      $@      "@      @      "@      @       @      �?       @                      �?      �?       @      �?                       @              @              @     �k@      4@     �k@      2@     @]@       @      X@              5@       @      4@      �?      @      �?      @                      �?      0@              �?      �?              �?      �?              Z@      0@      �?      @      �?      �?              �?      �?                      @     �Y@      (@     @X@       @      V@       @      S@              (@       @      @       @               @      @              "@              "@      @      @      @       @      @              @       @       @              �?       @      �?       @                      �?       @              @              @      @      �?      @      �?                      @      @                       @      3@     �T@              D@      3@     �E@      @      @      @                      @      (@     �C@      @     �A@      @       @               @      @               @     �@@      �?      ?@              ;@      �?      @      �?                      @      �?       @      �?      �?      �?                      �?              �?      @      @              @      @             �U@     �q@      5@     �f@      1@      X@      &@     @V@      @      1@      @      1@       @      @              @       @              @      &@      @      �?              �?      @                      $@       @              @      R@      @      K@             �E@      @      &@       @               @      &@              "@       @       @              �?       @      �?       @                      �?              2@      @      @      @              �?      @      �?      @      �?                      @              @      @     �U@             �P@      @      4@      @      3@      @       @      @                       @              1@      �?      �?      �?                      �?     @P@     �X@      O@     �N@      @      ,@              (@      @       @      @                       @      M@     �G@      I@      >@     �B@      @               @     �B@      @     �A@               @      @       @                      @      *@      9@      @      1@      @      @      �?      @              @      �?       @               @      �?               @                      (@      $@       @      @      @      @                      @      @      �?      @      �?       @               @      �?              �?       @              @               @      1@      @      @      @       @      @                       @              �?      @      ,@      @                      ,@      @     �B@       @      &@       @      �?              �?       @                      $@      �?      :@      �?       @      �?      @              @      �?       @               @      �?                      @              2@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKׅ�h~�B/         `                    �?U�ք�?�           ��@       ;                    @L@������?�            �r@       
                    I@ޗQ�~�?�            �i@                           @J@�q�q�?             (@              	          �����؇���X�?             @������������������������       �                     �?������������������������       �                     @       	                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?       8                   h@      �?             h@       '       	          ����?p�/E�f�?}            �g@                           �?�%IM��?c            �a@                           �?�E�����?=            �V@              
             �? �)���?8            @T@������������������������       �        4            �R@                            C@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@                          `]@@�0�!��?&            �I@                          `l@���Q��?             $@������������������������       �                     @                          �c@�q�q�?             @������������������������       �                     @                          p@�q�q�?             @������������������������       �                     �?                          `e@      �?              @������������������������       �                     �?������������������������       �                     �?       $                    �?,���i�?             �D@        !                   �q@�˹�m��?             C@������������������������       �                    �@@"       #                   �r@���Q��?             @������������������������       �                     @������������������������       �                      @%       &                     I@�q�q�?             @������������������������       �                      @������������������������       �                     �?(       7                    �?��|�5��?            �G@)       *       
             �?r�q��?             8@������������������������       �                     @+       ,       	          ����?b�2�tk�?             2@������������������������       �                     @-       2       	          ����?��S���?
             .@.       /                   �\@���Q��?             $@������������������������       �                     �?0       1                   �b@�q�q�?             "@������������������������       �                     @������������������������       �                     @3       6                    �E@z�G�z�?             @4       5                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        
             7@9       :                    d@      �?             @������������������������       �                     �?������������������������       �                     @<       G       
             �?�q�q��?:             X@=       >                    ]@؇���X�?            �A@������������������������       �                     �??       D                    �Q@�t����?             A@@       A       	            �? 7���B�?             ;@������������������������       �                     4@B       C       	          ����?؇���X�?             @������������������������       �                     �?������������������������       �                     @E       F                    �?և���X�?             @������������������������       �                     @������������������������       �                     @H       S                   �^@�'N��?&            �N@I       J                   `\@�FVQ&�?            �@@������������������������       �                     3@K       R                    �?؇���X�?	             ,@L       M                    �?���Q��?             @������������������������       �                     �?N       Q                   @^@      �?             @O       P                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@T       _                    �?���>4��?             <@U       ^       	          `ff@�ՙ/�?             5@V       ]                    @O@��Q��?             4@W       Z                    �?      �?
             ,@X       Y                   `k@      �?              @������������������������       �                      @������������������������       �                     @[       \                   �c@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @a       �                    �?Ƶ�pD�?            {@b       {       
             �?n60�F2�?r            �f@c       z                    `P@\`*�s�?5             U@d       i                    P@���5��?3            �S@e       h                   �_@؇���X�?             @f       g                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @j       k                   �b@�ӖF2��?-            �Q@������������������������       �                    �D@l       y                   �b@d��0u��?             >@m       x                    �?l��
I��?             ;@n       s                    �?��.k���?             1@o       p       	             �?r�q��?             @������������������������       �                     @q       r                   0l@      �?              @������������������������       �                     �?������������������������       �                     �?t       u                   `\@���|���?             &@������������������������       �                     @v       w                   �^@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     $@������������������������       �                     @������������������������       �                     @|       �                    �?n����W�?=            �X@}       ~       	          ����?,���i�?2            �T@������������������������       �                     E@       �                    ]@      �?             D@������������������������       �                     ,@�       �                     Q@�n_Y�K�?             :@�       �                   a@�q�q�?             8@�       �                     O@��.k���?             1@�       �                    c@�q�q�?	             (@������������������������       �                     @�       �                   �f@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   �[@z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   �`@ҳ�wY;�?             1@�       �                   �b@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                   0l@z�G�z�?             $@������������������������       �                     @�       �                   @n@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   P`@�uW��?�            `o@�       �                    Z@`<�Gf�?e             e@������������������������       �                     D@�       �                    �R@���f�?P             `@�       �       	          ����?      �?O             `@�       �       	          ����?8�Z$���?	             *@�       �                    @J@ףp=
�?             $@�       �                    _@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �^@�]���?F            �\@�       �                    �? >�֕�?            �A@�       �       
             �?�����?             5@������������������������       �                      @�       �                   Hs@�KM�]�?             3@�       �                   �h@�X�<ݺ?             2@������������������������       �                     (@�       �       	             �?r�q��?             @������������������������       �                      @�       �                    �K@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ,@������������������������       �        1             T@������������������������       �                     �?�       �       
             �?���?6            �T@�       �                   Pd@      �?             8@�       �                   `c@p�ݯ��?
             3@�       �                    �?�z�G��?             $@������������������������       �                     @�       �       	          033�?      �?             @������������������������       �                      @�       �                     N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@������������������������       �                     @�       �                   �U@\-��p�?(             M@������������������������       �                     @�       �       	          ����?�C��2(�?'            �K@�       �                   �n@PN��T'�?             ;@�       �                   �m@z�G�z�?             4@�       �                    �?�t����?
             1@�       �       	             �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     &@�       �                   �a@�q�q�?             @������������������������       �                     �?�       �                    @J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �Z@h�����?             <@�       �                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     9@�t�bh�h(h+K ��h-��R�(KK�KK��h_�Bp        t@     �y@     �k@      T@     �e@      ?@      @      @      �?      @      �?                      @      @      �?      @                      �?      e@      8@     �d@      5@     ``@      $@     @V@      �?      T@      �?     �R@              @      �?              �?      @              "@              E@      "@      @      @      @               @      @              @       @      �?      �?              �?      �?      �?                      �?      B@      @     �A@      @     �@@               @      @              @       @              �?       @               @      �?              B@      &@      *@      &@      @              @      &@              @      @       @      @      @              �?      @      @              @      @              �?      @      �?      �?              �?      �?                      @      7@              �?      @      �?                      @     �G@     �H@      >@      @              �?      >@      @      :@      �?      4@              @      �?              �?      @              @      @      @                      @      1@      F@       @      ?@              3@       @      (@       @      @      �?              �?      @      �?       @               @      �?                      �?              "@      .@      *@       @      *@      @      *@      @      @      @       @               @      @              �?      @              @      �?                      @      �?              @             �Y@     �t@     @S@     �Z@     �N@      7@     �N@      1@      �?      @      �?       @      �?                       @              @      N@      &@     �D@              3@      &@      3@       @      "@       @      @      �?      @              �?      �?              �?      �?              @      @              @      @       @      @                       @      $@                      @              @      0@     �T@      $@      R@              E@      $@      >@              ,@      $@      0@       @      0@       @      "@      @       @              @      @      �?      @                      �?      @      �?      �?      �?      �?                      �?      @                      @       @              @      &@      @      @      @                      @       @       @              @       @      @       @                      @      9@     @l@      @     �d@              D@      @      _@      @      _@       @      &@      �?      "@      �?      �?              �?      �?                       @      �?       @      �?                       @       @     @\@       @     �@@       @      3@               @       @      1@      �?      1@              (@      �?      @               @      �?      @              @      �?              �?                      ,@              T@      �?              4@      O@      (@      (@      @      (@      @      @      @              �?      @               @      �?      �?      �?                      �?              "@      @               @      I@      @              @      I@      @      7@      @      0@       @      .@       @      @              @       @                      &@       @      �?      �?              �?      �?      �?                      �?              @      �?      ;@      �?       @               @      �?                      9@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK�h~�B(5         �                    �?0����?�           ��@       Q       
             �?�ua��?           @{@       D                    �?��L��?�            �q@       #                    �?HP�s��?�            @o@                          �c@��-��ĳ?r            �e@       	                   @[@��	,UP�?A             W@                          �l@      �?             @������������������������       �                      @������������������������       �                      @
                           �?�zvܰ?>             V@                           @L@`Ql�R�?!            �G@������������������������       �                    �B@              	            �?ףp=
�?             $@������������������������       �                     @                          p`@�q�q�?             @������������������������       �                     �?������������������������       �                      @                          `a@������?            �D@������������������������       �                     @@                          `T@�<ݚ�?             "@������������������������       �                     �?                          �a@      �?              @              	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �?��Y��]�?1            �T@������������������������       �        &             Q@                           �?؇���X�?             ,@������������������������       �                     @       "                   �`@      �?              @        !                   �]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @$       -                    c@<�A+K&�?1             S@%       (                   @E@�����?             E@&       '       	          @33�?      �?             @������������������������       �                      @������������������������       �                      @)       *                    @M@�}�+r��?             C@������������������������       �                     6@+       ,                   @o@      �?
             0@������������������������       �                     ,@������������������������       �                      @.       C       	          ����?�������?             A@/       0                   �i@8^s]e�?             =@������������������������       �                      @1       >                    �?������?             ;@2       5                    ]@�q�q�?             2@3       4                    �?���Q��?             @������������������������       �                      @������������������������       �                     @6       =                   �b@�θ�?             *@7       8                    k@r�q��?             (@������������������������       �                     �?9       :                    �?�C��2(�?             &@������������������������       �                      @;       <                   Pf@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �??       @                    @M@�����H�?             "@������������������������       �                     @A       B                   @d@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @E       L                    �?�g�y��?             ?@F       K                   �b@r�q��?             2@G       J                     Q@�z�G��?             $@H       I                   �a@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @M       N                   �c@$�q-�?             *@������������������������       �                     @O       P                   �a@؇���X�?             @������������������������       �                     @������������������������       �                     �?R       ]       	          ����?n2�`���?b            `c@S       T                    �?�C��2(�?            �K@������������������������       �                    �F@U       X                    @F@      �?             $@V       W                   �d@      �?             @������������������������       �                     �?������������������������       �                     @Y       Z                   8p@�q�q�?             @������������������������       �                     @[       \                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?^       �                    �?Fx$(�?D             Y@_       �                   �t@���Q8�?5             T@`       �                   0o@      �?3             S@a       n                    �?^n����?'             N@b       e                    �F@"pc�
�?            �@@c       d                   �]@�q�q�?             @������������������������       �                     �?������������������������       �                      @f       g                   `k@�r����?             >@������������������������       �        	             1@h       i       	             �?�	j*D�?	             *@������������������������       �                      @j       m                    �?"pc�
�?             &@k       l                     J@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @o       ~                   �`@|��?���?             ;@p       w                   @l@�q�q�?
             .@q       v                   g@z�G�z�?             $@r       u                    �?      �?             @s       t                   @L@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @x       }                    `@���Q��?             @y       z                   �c@      �?             @������������������������       �                      @{       |       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?       �       	          ����?      �?	             (@������������������������       �                      @�       �                    �?ףp=
�?             $@�       �                    �?      �?             @�       �                    �P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     0@������������������������       �                     @�       �                    �?      �?             4@�       �                   @a@r�q��?             2@�       �       	          ����?��S�ۿ?             .@�       �                   `X@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                     P@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �       
             �?�q�� �?�            �r@�       �                   �b@�Q����?             D@�       �                    �?���Q��?            �A@������������������������       �                     @�       �                   Pj@      �?             <@�       �                    @L@؇���X�?             ,@������������������������       �                     @�       �                    �?      �?              @�       �                   �X@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                   �a@X�Cc�?
             ,@�       �                   �`@      �?              @�       �       	          033�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   `_@r�q��?             @������������������������       �                     @�       �                   @b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?�����?�             p@�       �                    �?������?            �F@�       �                    �E@� �	��?             9@������������������������       �                     @�       �       	             �?�z�G��?             4@�       �       	             �?X�<ݚ�?             "@������������������������       �                     �?�       �                    �J@      �?              @������������������������       �                      @�       �                    �?r�q��?             @�       �                   @_@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �`@�C��2(�?             &@������������������������       �                      @�       �                    �?�q�q�?             @�       �                    @H@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    c@P���Q�?             4@������������������������       �                     3@������������������������       �                     �?�       �                   �b@�����?�            �j@�       �                    �?��S�ۿ?�            @j@�       �                   �Z@,_ʯ08�?b            �c@������������������������       �                      @�       �                    \@�E����?a            �c@�       �                   `[@X�EQ]N�?            �E@�       �                   �W@Pa�	�?            �@@������������������������       �        	             0@�       �                   @X@�IєX�?             1@�       �                    �?z�G�z�?             @������������������������       �                      @�       �                   (q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             (@�       �                   �k@���Q��?             $@������������������������       �                     @�       �       	          ����?և���X�?             @������������������������       �                      @�       �                    �K@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   0f@�}�+r��?E            �\@������������������������       �                     9@�       �       	          ����?���M�?5            @V@�       �                   �`@�p ��?            �D@�       �                    �?�����?             3@�       �                   �m@z�G�z�?             .@�       �                   �l@      �?              @�       �                    �I@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �a@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     6@������������������������       �                     H@�       �                   s@���J��?!            �I@������������������������       �                     F@�       �                    �P@؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK�KK��h_�B0        u@     �x@     r@     `b@     �n@     �A@     �l@      4@     �d@      @     �U@      @       @       @       @                       @     @U@      @      G@      �?     �B@              "@      �?      @               @      �?              �?       @             �C@       @      @@              @       @              �?      @      �?      �?      �?              �?      �?              @              T@       @      Q@              (@       @      @              @       @      �?       @      �?                       @      @             �O@      *@      C@      @       @       @       @                       @      B@       @      6@              ,@       @      ,@                       @      9@      "@      4@      "@               @      4@      @      (@      @       @      @       @                      @      $@      @      $@       @              �?      $@      �?       @               @      �?              �?       @                      �?       @      �?      @               @      �?              �?       @              @              0@      .@      .@      @      @      @      @      �?      @                      �?               @       @              �?      (@              @      �?      @              @      �?             �E@      \@      @      I@             �F@      @      @      @      �?              �?      @               @      @              @       @      �?       @                      �?      C@      O@      7@     �L@      3@     �L@      3@     �D@      @      ;@       @      �?              �?       @              @      :@              1@      @      "@       @               @      "@       @      @              @       @                      @      *@      ,@      $@      @       @       @       @       @      �?       @      �?                       @      �?              @               @      @      �?      @               @      �?      �?      �?                      �?      �?              @      "@       @              �?      "@      �?      @      �?      �?              �?      �?                       @              @              0@      @              .@      @      .@      @      ,@      �?      @      �?              �?      @               @              �?       @               @      �?                       @     �G@     `o@      3@      5@      ,@      5@      @              @      5@       @      (@              @       @      @       @       @               @       @                      @      @      "@      @      @      �?      @              @      �?              @              �?      @              @      �?      �?              �?      �?              @              <@     �l@      (@     �@@      &@      ,@      @              @      ,@      @      @              �?      @      @               @      @      �?      @      �?              �?      @               @              �?      $@               @      �?       @      �?      �?              �?      �?                      �?      �?      3@              3@      �?              0@     �h@      ,@     �h@      *@     @b@       @              &@     @b@      @      C@      �?      @@              0@      �?      0@      �?      @               @      �?       @      �?                       @              (@      @      @              @      @      @       @               @      @       @                      @      @      [@              9@      @     �T@      @     �A@      @      *@      @      (@      @      @      �?      @              @      �?               @                      @      @      �?      @                      �?              6@              H@      �?      I@              F@      �?      @              @      �?               @      �?       @                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKŅ�h~�B+         N                    �?�+	G�?�           ��@              
             �?�@o-4�?�            �s@                          �g@P���Q�?y             i@                          �O@��:x�ٳ?x            �h@������������������������       �                     @                          �a@`�E���?u            @h@������������������������       �        %             O@                          �a@Pa�	�?P            �`@	       
                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �? g�yB�?N             `@                           �?�x�E~�?8            @V@������������������������       �                    �E@                          �e@�nkK�?             G@                          @[@      �?             @@                          @Y@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?(;L]n�?             >@                          �e@���7�?             6@������������������������       �                     3@                            H@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     ,@������������������������       �                     D@������������������������       �                      @       C                    �?�>4ևF�?G             \@       *                    @K@�c�Α�?8            �U@        )                    �?l��[B��?             =@!       &                    �?r�q��?             2@"       %                    �D@����X�?             @#       $                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @'       (                     F@�C��2(�?
             &@������������������������       �                     �?������������������������       �        	             $@������������������������       �                     &@+       6                    �?д>��C�?#             M@,       3                   �a@�X����?             6@-       2                   P`@��S�ۿ?
             .@.       /                   �p@z�G�z�?             @������������������������       �                     @0       1                   @[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@4       5                    �K@؇���X�?             @������������������������       �                     �?������������������������       �                     @7       >                   @L@�8��8��?             B@8       =                    �?���Q��?             @9       :                    ]@�q�q�?             @������������������������       �                     �?;       <                    �P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @?       @                    c@�g�y��?             ?@������������������������       �                     5@A       B                    [@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@D       M                    �?�+e�X�?             9@E       L                    �?�q�q�?             8@F       G                   �Z@�㙢�c�?             7@������������������������       �                     @H       K                   �g@P���Q�?             4@I       J       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             2@������������������������       �                     �?������������������������       �                     �?O       �                    �?.�����?           `z@P       w       	          ����?�+Ze��?�            �u@Q       r                    �?�D#���?K            �\@R       k       
             �?X�<ݚ�?7            @T@S       T                   `X@����X�?             E@������������������������       �                     @U       ^                    c@�θ�?            �C@V       [                    �?ȵHPS!�?             :@W       X                    �?���N8�?             5@������������������������       �        	             ,@Y       Z                    T@؇���X�?             @������������������������       �                     �?������������������������       �                     @\       ]                    �?���Q��?             @������������������������       �                      @������������������������       �                     @_       j                    b@��
ц��?
             *@`       a                    �A@���|���?             &@������������������������       �                     �?b       e                    �?�z�G��?             $@c       d                   `Z@؇���X�?             @������������������������       �                     �?������������������������       �                     @f       i       	          @33�?�q�q�?             @g       h                   �e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @l       o                    �O@8�Z$���?            �C@m       n       	          ����?      �?             @@������������������������       �                     ?@������������������������       �                     �?p       q                   �j@����X�?             @������������������������       �                      @������������������������       �                     @s       t                   �b@l��\��?             A@������������������������       �                     <@u       v                   �c@      �?             @������������������������       �                     @������������������������       �                     @x       �                   �c@��i���?�            �l@y       �       
             �?$Nz�{�?�             k@z       {                    �H@      �?             (@������������������������       �                     @|       }                   �\@�q�q�?             "@������������������������       �                     �?~                           �?      �?              @������������������������       �                     @������������������������       �                      @�       �                    �?�À���?�            �i@�       �                    �R@ȑ����?N            @]@�       �                    �L@ �^�@̩?M             ]@������������������������       �        3            �S@�       �                   q@�˹�m��?             C@������������������������       �                     >@�       �                   �a@      �?              @�       �                   �S@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �                   0a@`���i��?9             V@�       �                    @O@hA� �?0            �Q@�       �       	          `ff@���J��?"            �I@������������������������       �                    �D@�       �                   �\@ףp=
�?             $@�       �                   �[@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �O@�KM�]�?             3@�       �                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     0@�       �                    �H@�<ݚ�?	             2@������������������������       �                     @������������������������       �                     ,@�       �                   �_@X�Cc�?             ,@������������������������       �                     @�       �                   `a@      �?             $@������������������������       �                     @�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �       
             �?p�ݯ��?.             S@�       �                   �^@�J�4�?             9@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @�       �       	             �?�}�+r��?             3@�       �                   �b@�IєX�?	             1@������������������������       �                     $@�       �                    �N@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?L紂P�?            �I@�       �                   (s@$G$n��?            �B@�       �       	          `ff@l��\��?             A@�       �                     Q@�FVQ&�?            �@@�       �                    �?      �?             @@�       �                   �X@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     8@������������������������       �                     �?������������������������       �                     �?�       �       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	          ����?؇���X�?
             ,@�       �                   `@����X�?             @������������������������       �                     @�       �                   8p@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�BP       `t@     �y@      m@     �S@     �g@      $@     �g@       @              @     �g@      @      O@              `@      @      �?       @               @      �?             �_@       @     �U@       @     �E@              F@       @      >@       @      �?      �?      �?                      �?      =@      �?      5@      �?      3@               @      �?       @                      �?       @              ,@              D@                       @     �E@     @Q@      8@     �O@      ,@      .@      @      .@       @      @       @       @               @       @                      @      �?      $@      �?                      $@      &@              $@      H@      @      .@      �?      ,@      �?      @              @      �?      �?              �?      �?                      $@      @      �?              �?      @              @     �@@       @      @       @      �?      �?              �?      �?      �?                      �?               @      �?      >@              5@      �?      "@      �?                      "@      3@      @      3@      @      3@      @              @      3@      �?      �?      �?      �?                      �?      2@                      �?              �?     @W@     �t@     @P@     �q@     �C@      S@      B@     �F@      >@      (@              @      >@      "@      7@      @      4@      �?      ,@              @      �?              �?      @              @       @               @      @              @      @      @      @              �?      @      @      @      �?              �?      @              �?       @      �?      �?              �?      �?                      �?               @      @     �@@      �?      ?@              ?@      �?              @       @               @      @              @      ?@              <@      @      @      @                      @      :@     �i@      1@      i@      @      @              @      @      @              �?      @       @      @                       @      &@     @h@      @     @\@      @     @\@             �S@      @     �A@              >@      @      @      �?      @      �?                      @       @              �?              @     @T@      @     �P@      �?      I@             �D@      �?      "@      �?       @               @      �?                      @       @      1@       @      �?       @                      �?              0@      @      ,@      @                      ,@      "@      @      @              @      @              @      @      �?      @                      �?      <@      H@      5@      @      @      @      @                      @      2@      �?      0@      �?      $@              @      �?              �?      @               @              @      F@      @      @@      @      ?@       @      ?@      �?      ?@      �?      @              @      �?                      8@      �?              �?               @      �?       @                      �?       @      (@       @      @              @       @       @               @       @                      @�t�bub��(     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKӅ�h~�B(.         |                    �?6������?�           ��@       [       	          ����?�C�"��?"           �{@                          `_@n(��"�?�            v@                           �?��
ц��?.            @P@                           @K@      �?$             H@              
             �?r�q��?             8@       
                    �?$�q-�?             *@       	       	             �?ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     @                           �?�C��2(�?             &@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@                          8w@�q�q�?             8@                           Z@�㙢�c�?             7@              
             �?      �?              @������������������������       �                     @������������������������       �                     @              
             �?��S�ۿ?	             .@                          @\@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@������������������������       �                     �?������������������������       �        
             1@       D       
             �?F��ӭ��?�             r@       /                    �?     ��?�             l@       .                    f@!�;��?p            �e@        -                   �c@��˼��?o             e@!       ,                    �?���N8�?8             U@"       +                   �c@@4և���?$             L@#       *                    �?�O4R���?#            �J@$       %                   �a@h�����?             <@������������������������       �        	             ,@&       '                     L@@4և���?             ,@������������������������       �        	             &@(       )                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     9@������������������������       �                     @������������������������       �                     <@������������������������       �        7            @U@������������������������       �                     @0       1                   Pe@R�}e�.�?              J@������������������������       �                     $@2       ?                     L@�q�q�?             E@3       <       	          433�?�������?             >@4       ;                    @F@d}h���?             <@5       :                   �b@ҳ�wY;�?	             1@6       9                    ]@������?             .@7       8                    �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �        	             &@=       >                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?@       C                    �?�q�q�?             (@A       B                   �j@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @E       F                   �f@     ��?&             P@������������������������       �        	             1@G       R                    �?��V�I��?            �G@H       I                    �?8�A�0��?             6@������������������������       �                     @J       Q                   �d@     ��?             0@K       P                    �L@�q�q�?             "@L       M       	          ����?؇���X�?             @������������������������       �                     @N       O                   ``@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @S       Z                    �N@`�Q��?             9@T       U       	          ����?      �?
             0@������������������������       �                     @V       Y       	          ����?z�G�z�?             $@W       X                    �K@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     "@\       o                   �c@���?>            @V@]       l                    �?�k�'7��?(            �L@^       a                   pe@��R[s�?            �A@_       `                    `@����X�?             @������������������������       �                     @������������������������       �                      @b       g                    �?؇���X�?             <@c       d                   �^@      �?              @������������������������       �                     @e       f       	             @���Q��?             @������������������������       �                     @������������������������       �                      @h       i                     P@P���Q�?             4@������������������������       �                     2@j       k                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?m       n                   �b@���7�?             6@������������������������       �                     5@������������������������       �                     �?p       {       	             @     ��?             @@q       t                    �?�q�q�?             8@r       s                   �e@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?u       z                    e@և���X�?	             ,@v       y                    �?���!pc�?             &@w       x                    �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @}       �                    �?v���a�?�            @r@~       �                    �?X�<ݚ�?             2@       �                   �c@"pc�
�?             &@�       �                   �`@ףp=
�?             $@�       �                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    d@؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?d/�@7�?�             q@�       �                   �b@pTjD��?�             n@�       �       
             �?��g�?�            @k@�       �                   (r@     ��?             0@�       �       	          ����?�q�q�?
             (@������������������������       �                     @�       �                    �?�<ݚ�?             "@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �U@��^M}�?�            @i@������������������������       �                      @�       �                   Xs@`2U0*��?�             i@�       �                    �K@P�p�_�?w            `f@�       �                   �l@ ��WV�?2            �S@������������������������       �                     G@�       �                   �l@     ��?             @@������������������������       �                     �?�       �                    �?`Jj��?             ?@������������������������       �                     1@�       �                   �`@؇���X�?	             ,@�       �       	          ���@�8��8��?             (@������������������������       �                     $@�       �                    �J@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �F@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          hff�?�����?E            @Y@�       �       	          ����?@4և���?
             ,@������������������������       �        	             *@������������������������       �                     �?������������������������       �        ;            �U@�       �                    �?��s����?             5@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �R@�IєX�?             1@������������������������       �        
             0@������������������������       �                     �?�       �                    �C@\X��t�?             7@������������������������       �                     @�       �                    _@�\��N��?             3@������������������������       �                     @�       �                   �g@     ��?	             0@������������������������       �                     @�       �                   �i@��
ц��?             *@�       �                   @`@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   �c@����X�?             @������������������������       �                      @������������������������       �                     @�       �                    �?�q�q�?            �@@�       �                    �H@
j*D>�?             :@�       �                    �?�<ݚ�?             "@�       �                   �`@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                   �`@������?             1@�       �       	          @33�?���|���?             &@������������������������       �                     @�       �                   @_@      �?              @������������������������       �                      @�       �       
             �?�q�q�?             @������������������������       �                     �?�       �                   h@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B0       �t@     �x@     0r@     �b@     �p@     @V@     �A@      >@      2@      >@      *@      &@      (@      �?      "@      �?      "@                      �?      @              �?      $@      �?      �?              �?      �?                      "@      @      3@      @      3@      @      @      @                      @      �?      ,@      �?       @               @      �?                      (@      �?              1@             �l@     �M@     `i@      5@     �d@      @     �d@      @      T@      @      J@      @      J@      �?      ;@      �?      ,@              *@      �?      &@               @      �?              �?       @              9@                      @      <@             @U@                      @      C@      ,@      $@              <@      ,@      7@      @      6@      @      &@      @      &@      @      @      @      @                      @      @                       @      &@              �?      �?      �?                      �?      @      @      @       @               @      @                      @      :@      C@              1@      :@      5@      "@      *@      @              @      *@      @      @      �?      @              @      �?      �?      �?                      �?       @                      @      1@       @       @       @              @       @       @      @       @      @                       @      @              "@              ;@      O@      $@     �G@      "@      :@      @       @      @                       @      @      8@      @      @              @      @       @      @                       @      �?      3@              2@      �?      �?      �?                      �?      �?      5@              5@      �?              1@      .@      1@      @      "@      �?      "@                      �?       @      @       @      @      @      @              @      @              @                      @               @      F@      o@       @      $@       @      "@      �?      "@      �?       @               @      �?                      @      �?              @      �?      @                      �?      B@     �m@      9@      k@      .@     `i@      @      &@      @      @      @               @      @       @       @       @                       @              @              @      $@      h@       @               @      h@      @     �e@      @     �R@              G@      @      =@      �?               @      =@              1@       @      (@      �?      &@              $@      �?      �?      �?                      �?      �?      �?              �?      �?              �?      Y@      �?      *@              *@      �?                     �U@      @      1@      @      �?      @                      �?      �?      0@              0@      �?              $@      *@              @      $@      "@      @              @      "@              @      @      @      @      �?              �?      @               @      @       @                      @      &@      6@      &@      .@      @       @      @       @               @      @               @              @      *@      @      @              @      @      @       @               @      @      �?              �?      @      �?                      @              @              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJQY%hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK߅�h~�B�0         �                    �?�Z���?�           ��@       C                    �?~�Q7:�?           �z@       $       
             �?�d���?�             n@              	            �?p�u$v��?u            �f@                           �?PL��V�?a            �b@                           �?�H�I���?J            @\@������������������������       �        -            �Q@                          @[@�Ń��̧?             E@	       
                    �J@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                    �C@                          pg@ >�֕�?            �A@                          `c@г�wY;�?             A@������������������������       �                     @@                          �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                           U@�'�`d�?            �@@������������������������       �                      @       #                    �?�חF�P�?             ?@                           �?�GN�z�?             6@                          @b@����X�?             ,@                            K@�q�q�?             @������������������������       �                     �?                          p`@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @                            �?      �?              @������������������������       �                     @!       "                    a@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@%       >                    �?����*��?'            �M@&       /                    �F@P����?             C@'       .                    �?X�<ݚ�?             "@(       -                   �_@�q�q�?             @)       ,                   �b@z�G�z�?             @*       +                    �C@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @0       1                     J@�c�Α�?             =@������������������������       �                     @2       7                    �?�LQ�1	�?             7@3       6                    �?���Q��?             $@4       5                   �^@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @8       =                   xp@�	j*D�?
             *@9       :                   �b@      �?	             (@������������������������       �                     @;       <                   �_@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �??       B                    �H@�����?             5@@       A                    b@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �        	             0@D       q                    �?,�[I'��?w            �g@E       b       
             �?<ݚ)�?^             b@F       a                   �b@���Q��?*            @P@G       ^       	            �?�-ῃ�?(            �N@H       O                   @E@�D��?             �H@I       N                   �_@z�G�z�?             $@J       K                   �X@�q�q�?             @������������������������       �                     @L       M       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @P       ]       	          ����?�ݜ�?            �C@Q       R                   �b@д>��C�?             =@������������������������       �        
             ,@S       X                   �d@�q�q�?             .@T       U                    @H@և���X�?             @������������������������       �                      @V       W                    b@���Q��?             @������������������������       �                     @������������������������       �                      @Y       \                   f@      �?              @Z       [                   Pe@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@_       `                   �a@      �?             (@������������������������       �                     "@������������������������       �                     @������������������������       �                     @c       n                   �d@86��Z�?4            �S@d       e       	             �?xL��N�?1            �R@������������������������       �                     D@f       m                   a@l��\��?             A@g       l                   @v@�S����?             3@h       i                   pc@�����H�?             2@������������������������       �                     .@j       k                    X@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �        
             .@o       p       	          ����?���Q��?             @������������������������       �                     @������������������������       �                      @r                          �c@�X����?             F@s       ~                    �?|��?���?             ;@t       u       
             �?8�A�0��?             6@������������������������       �                     @v       }                    `P@���Q��?
             .@w       x                   �Z@"pc�
�?             &@������������������������       �                     �?y       z                   �c@ףp=
�?             $@������������������������       �                      @{       |                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     1@�       �                   �b@$��n�?�             s@�       �                    �?؇���X�?�            q@�       �       	          433�?      �?	             (@�       �       
             �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                     K@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�=C|F�?�            Pp@�       �                    �?�h��?|            �g@�       �                    @N@�+ت�M�?k            �c@�       �                    [@�8�So��?Q            @^@������������������������       �                     @�       �                   �e@�y��*�?N             ]@�       �       
             �?hdpZ�L�?L            @\@�       �       	          ����?և���X�?             @������������������������       �                     @�       �                   �\@      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �h@��-#���?F            �Z@������������������������       �                    �D@�       �       	          ����?��ɉ�?-            @P@�       �                    l@�z�G��?             4@�       �       	             �?�C��2(�?             &@������������������������       �                     "@�       �                    �I@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �J@X�<ݚ�?             "@�       �                   �`@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   j@��S�ۿ?!            �F@������������������������       �                     �?�       �       	          033@���7�?              F@������������������������       �                    �A@�       �                   8p@�<ݚ�?             "@������������������������       �                     @�       �                    �J@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   Xp@�?�|�?            �B@������������������������       �                     :@�       �                   �p@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@�       �       	          433�?f���M�?             ?@������������������������       �                     @�       �                   �`@� �	��?             9@�       �                    @H@�	j*D�?             *@������������������������       �                      @�       �                   h@"pc�
�?             &@������������������������       �                     @�       �                    _@����X�?             @������������������������       �                     @�       �                   @_@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �H@r�q��?             (@�       �                   �]@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                    �R@������?-             R@�       �       
             �? ��PUp�?,            �Q@�       �                   �^@z�G�z�?             @������������������������       �                     @�       �                   �r@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        (            �P@������������������������       �                     �?�       �                   `c@�q�q�?            �@@�       �                    b@�8��8��?             (@������������������������       �                     @�       �                   �q@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�G��l��?             5@�       �                   `d@X�Cc�?             ,@������������������������       �                      @�       �                   �q@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�        u@     �x@     Pq@     �b@     `i@     �B@     `e@      $@      b@      @      \@      �?     �Q@             �D@      �?       @      �?              �?       @             �C@             �@@       @     �@@      �?      @@              �?      �?              �?      �?                      �?      :@      @               @      :@      @      1@      @      $@      @       @      @      �?              �?      @              @      �?               @              @      �?      @              @      �?              �?      @              "@              @@      ;@      *@      9@      @      @       @      @      �?      @      �?      �?              �?      �?                      @      �?              @               @      5@              @       @      .@      @      @      @      @              @      @                       @      @      "@      @      "@              @      @       @               @      @              �?              3@       @      @       @      @                       @      0@             �R@     �\@      F@      Y@     �C@      :@     �C@      6@      B@      *@       @       @       @      @              @       @      �?       @                      �?              @      A@      @      8@      @      ,@              $@      @      @      @               @      @       @      @                       @      @      �?      @      �?      @                      �?      @              $@              @      "@              "@      @                      @      @     �R@      @     �Q@              D@      @      ?@      @      0@       @      0@              .@       @      �?              �?       @              �?                      .@       @      @              @       @              >@      ,@      *@      ,@      *@      "@      @              @      "@       @      "@      �?              �?      "@               @      �?      �?              �?      �?              @                      @      1@             �N@     �n@     �C@     @m@      @      @      @      �?      @                      �?      �?      @      �?                      @     �@@     �l@      ?@     �c@      4@     @a@      3@     �Y@      @              ,@     �Y@      (@     @Y@      @      @              @      @      �?       @              �?      �?      �?                      �?      "@     @X@             �D@      "@      L@      @      ,@      �?      $@              "@      �?      �?              �?      �?              @      @      @      @              @      @               @              @      E@      �?               @      E@             �A@       @      @              @       @       @       @                       @       @      �?       @                      �?      �?      B@              :@      �?      $@      �?                      $@      &@      4@              @      &@      ,@      "@      @               @      "@       @      @              @       @      @              �?       @      �?                       @       @      $@       @       @               @       @                       @       @     �Q@      �?     �Q@      �?      @              @      �?      �?      �?                      �?             �P@      �?              6@      &@      &@      �?      @              @      �?              �?      @              &@      $@      @      "@               @      @      �?      @                      �?      @      �?      @                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��fbhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKυ�h~�BH-         L                    �?�#i����?�           ��@              
             �?�� ~E��?�            s@       
                    I@�8��8��?y            �i@                           ^@8�Z$���?             *@������������������������       �                     �?                          Pb@�8��8��?             (@������������������������       �                     "@       	                    �J@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           @L@�w��3(�?s            �g@                          @[@���=��?]            �b@                           �?�C��2(�?             &@������������������������       �                     @                          �Z@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �        X            `a@              	          833@,���i�?            �D@                          p@$�q-�?            �C@������������������������       �                     7@                          �c@     ��?	             0@                          @a@�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @       =                    �?:�o���?@            @Y@                          �Z@      �?&             L@������������������������       �                     @       (                   ph@r�z-��?$            �J@        !       	          @33�?��S���?	             .@������������������������       �                      @"       '                   d@��
ц��?             *@#       $                    �?      �?              @������������������������       �                     @%       &                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @)       *                   �[@�d�����?             C@������������������������       �                     @+       ,                   �j@z�G�z�?            �A@������������������������       �                     &@-       <       	          ��� @�q�q�?             8@.       3       	          ����?��s����?             5@/       0                   @b@���Q��?             @������������������������       �                     �?1       2                     H@      �?             @������������������������       �                     �?������������������������       �                     @4       5                    _@      �?             0@������������������������       �                     �?6       7                    �L@��S�ۿ?             .@������������������������       �        	             &@8       ;                   �z@      �?             @9       :                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @>       K                   �b@������?            �F@?       F                   �`@�?�'�@�?             C@@       E                   P`@ ��WV�?             :@A       B                   �_@�8��8��?             (@������������������������       �                     @C       D       	             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             ,@G       H                     M@�q�q�?             (@������������������������       �                     @I       J                    �?և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @M       �       	          ����?�f|��?           �z@N       {       
             �?      �?f            �c@O       f                    �L@�?�Ʋ(�?8            @W@P       e                    �?     8�?%             P@Q       `                    @F@F�4�Dj�?"            �M@R       S                    T@�n_Y�K�?             :@������������������������       �                     @T       U                   pb@���N8�?             5@������������������������       �                     @V       _                    �?�q�q�?             .@W       \                    ]@�n_Y�K�?	             *@X       Y                   �c@z�G�z�?             @������������������������       �                     @Z       [                    �E@      �?              @������������������������       �                     �?������������������������       �                     �?]       ^                   �b@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @a       b                   �d@Pa�	�?            �@@������������������������       �                     >@c       d                   �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @g       v       	          833�?l��[B��?             =@h       s                   �b@��Q��?             4@i       l                    _@      �?
             0@j       k       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?m       n                   @Z@8�Z$���?             *@������������������������       �                     �?o       r                    �M@�8��8��?             (@p       q                   f@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @t       u                   `^@      �?             @������������������������       �                     @������������������������       �                     �?w       x                    �?�����H�?             "@������������������������       �                     @y       z                   �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @|       �       	          ����?�z����?.            @P@}       ~                    �?@�E�x�?$            �H@������������������������       �                    �E@       �                   `^@r�q��?             @������������������������       �                     @�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �_@      �?
             0@������������������������       �                     @�       �       	          ����?r�q��?             (@�       �                    �?�q�q�?             @�       �                    X@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �c@,7���v�?�            �p@�       �                    �?���>�?�            �n@�       �                    �?X'"7��?�             k@�       �                   pj@D��*�4�?c            @a@�       �                    \@���@��?            �B@�       �                    �F@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    @L@      �?             @@������������������������       �        	             *@�       �       
             �?���y4F�?             3@�       �                   �\@      �?             @������������������������       �                     �?�       �       	          033�?�q�q�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�r����?             .@������������������������       �                     �?�       �                    �?@4և���?             ,@������������������������       �                      @�       �                   �`@r�q��?             @�       �                   @_@      �?             @������������������������       �                     �?�       �                    �L@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   �v@��:�-�?D            @Y@�       �                   `a@`�LVXz�?B            �X@������������������������       �        2            @S@�       �                   �[@���7�?             6@�       �                   �a@�q�q�?             @�       �                    @K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     3@�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        -            �S@�       �                    �P@�z�G��?             >@�       �                   �`@���B���?             :@�       �                   @_@���|���?             &@������������������������       �                     @������������������������       �                     @�       �                    �H@��S�ۿ?             .@�       �                   �k@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             *@������������������������       �                     @�       �                   `T@���Q��?             9@������������������������       �                     @�       �                   �o@X�<ݚ�?             2@�       �                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @�       �                    b@      �?              @�       �                   �c@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       `u@     �x@     @m@     �Q@     `g@      1@       @      &@      �?              �?      &@              "@      �?       @               @      �?              g@      @     �b@      �?      $@      �?      @              @      �?      @                      �?     `a@              B@      @      B@      @      7@              *@      @      @      @      @                      @      @                       @     �G@      K@     �A@      5@              @     �A@      2@      @       @               @      @      @      @      �?      @              �?      �?              �?      �?                      @      <@      $@              @      <@      @      &@              1@      @      1@      @      @       @              �?      @      �?              �?      @              ,@       @              �?      ,@      �?      &@              @      �?      �?      �?              �?      �?               @                      @      (@     �@@      @     �@@      �?      9@      �?      &@              @      �?      @              @      �?                      ,@      @       @              @      @      @      @                      @      @              [@     t@     �S@     �S@      Q@      9@     �J@      &@      H@      &@      0@      $@              @      0@      @      @              $@      @       @      @      �?      @              @      �?      �?      �?                      �?      @      �?      @                      �?       @              @@      �?      >@               @      �?       @                      �?      @              .@      ,@      @      *@      @      (@       @      �?       @                      �?       @      &@      �?              �?      &@      �?      @              @      �?                       @      @      �?      @                      �?       @      �?      @               @      �?              �?       @              &@      K@      �?      H@             �E@      �?      @              @      �?      �?      �?                      �?      $@      @              @      $@       @      @       @      @      �?              �?      @                      �?      @              =@     @n@      3@     `l@      $@     �i@      $@      `@       @      =@      @      �?              �?      @              @      <@              *@      @      .@       @       @              �?       @      �?      �?              �?      �?      �?                      �?       @      *@      �?              �?      *@               @      �?      @      �?      @              �?      �?       @      �?                       @               @       @     �X@      �?     �X@             @S@      �?      5@      �?       @      �?      �?      �?                      �?              �?              3@      �?      �?      �?                      �?             �S@      "@      5@      @      5@      @      @      @                      @      �?      ,@      �?      �?              �?      �?                      *@      @              $@      .@              @      $@       @       @       @       @                       @       @      @      �?      @      �?                      @      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ$�phG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKυ�h~�BH-         X       
             �?"��G,�?�           ��@       E                    �?DE��2{�?�            �r@                           �?6C�d�?�            �o@              	             @Pq�����?m            @e@                          �g@�|�%T�?l             e@                           �?h�����?k             e@              	            �? �h�7W�?C            �Z@                          @[@`Ӹ����?9            �V@	       
                   �Z@�q�q�?             "@������������������������       �                     @������������������������       �                     @                          �t@ �)���?5            @T@������������������������       �        4             T@������������������������       �                     �?                          @a@      �?
             0@������������������������       �                      @                          @b@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �        (             O@������������������������       �                     �?������������������������       �                     �?       *                   �j@��]�T��?2            �T@       '                    i@�eP*L��?            �@@       &                    �?�q�q�?             8@                           �?�G��l��?             5@                           @L@ףp=
�?             $@������������������������       �                     @                           �M@�q�q�?             @������������������������       �                     �?������������������������       �                      @        !                    �H@"pc�
�?             &@������������������������       �                     @"       #                   @Z@���Q��?             @������������������������       �                      @$       %                     P@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @(       )                    _@�����H�?             "@������������������������       �                     �?������������������������       �                      @+       >                   �b@ \� ���?            �H@,       ;                    �?�T|n�q�?            �E@-       8                    �O@�KM�]�?             C@.       /                    �?`Jj��?             ?@������������������������       �                     $@0       1                    @F@�����?             5@������������������������       �                     �?2       3                   �^@P���Q�?
             4@������������������������       �                     &@4       5                   �d@�����H�?             "@������������������������       �                     @6       7                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?9       :                   Pc@����X�?             @������������������������       �                     @������������������������       �                      @<       =       	          ����?���Q��?             @������������������������       �                      @������������������������       �                     @?       D                    �?r�q��?             @@       A                    �?z�G�z�?             @������������������������       �                      @B       C                   �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?F       I                    �?r�q��?             H@G       H                    V@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@J       S                    �?P����?             C@K       R                   ``@�n_Y�K�?             :@L       Q                    _@���!pc�?
             6@M       P                    �J@ҳ�wY;�?             1@N       O                     F@�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @T       W                    `P@      �?             (@U       V       	          ����?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                      @Y       h                    �?�*�@P��?            {@Z       c                    @L@l��[B��?             =@[       b                    �?�q�q�?             5@\       a                   Pl@��
ц��?	             *@]       `                    Y@؇���X�?             @^       _                   �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @d       g                   P`@      �?              @e       f                   Po@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @i       �                    �?T&ss��?�            Py@j       �                   �a@���	D�?�            �u@k       �                   @d@H�te�?�            `q@l       o                   �Q@�5ĉ*�?�            `o@m       n                    �?���Q��?             @������������������������       �                      @������������������������       �                     @p       �                    �?0��P�?�            �n@q       r                   �h@$�q-�?P            @`@������������������������       �                     �H@s       t                   @i@�$�����?0            @T@������������������������       �                     @u       v                    @K@�:�^���?/            �S@������������������������       �                     ?@w       �                   �[@��0{9�?            �G@x       {                    �K@��+7��?             7@y       z       	             �?�q�q�?             @������������������������       �                     @������������������������       �                      @|       }                   �Y@�t����?             1@������������������������       �                     &@~                          �`@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   �`@ �q�q�?             8@������������������������       �                     3@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    m@���"�?C             ]@�       �                   �\@�k~X��?*             R@�       �                    �?�IєX�?             1@�       �                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@������������������������       �                    �K@�       �                   �m@�C��2(�?             F@������������������������       �                      @�       �                    �J@���N8�?             E@�       �                    @J@z�G�z�?             $@������������������������       �                     @�       �                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @@������������������������       �                     ;@�       �                    �K@�q�q�?(             R@�       �                   �i@�IєX�?             A@������������������������       �        	             ,@�       �                    �?ףp=
�?
             4@�       �                   �m@z�G�z�?             @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �Z@��S�ۿ?             .@������������������������       �                     �?������������������������       �                     ,@�       �                   �`@P����?             C@�       �                   Pb@D�n�3�?
             3@������������������������       �                     @�       �                    �?�n_Y�K�?             *@�       �       	          033�?�q�q�?             (@������������������������       �                     @�       �                   pj@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                    �M@�KM�]�?             3@�       �       	          433�?�q�q�?             @������������������������       �                     �?�       �                    c@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@�       �                   `c@�eP*L��?&            �K@�       �                   �c@X�<ݚ�?!            �F@�       �                    `P@      �?             D@�       �       	          ����?      �?             @@�       �       	          833�?��
ц��?             :@�       �                    �?      �?              @�       �                   @n@z�G�z�?             @������������������������       �                     @�       �                   @b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �[@b�2�tk�?             2@������������������������       �                     �?�       �                   `X@ҳ�wY;�?             1@������������������������       �                     �?�       �                   �q@     ��?
             0@�       �                   �^@�eP*L��?             &@������������������������       �                      @�       �                    @M@�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       @s@     �z@     �m@      P@     �j@      C@     @d@       @     @d@      @     @d@      @      Y@      @     �U@      @      @      @      @                      @      T@      �?      T@                      �?      ,@       @       @              @       @               @      @              O@                      �?              �?      J@      >@      .@      2@      ,@      $@      &@      $@      "@      �?      @               @      �?              �?       @               @      "@              @       @      @               @       @      �?       @                      �?      @              �?       @      �?                       @     �B@      (@      B@      @      A@      @      =@       @      $@              3@       @              �?      3@      �?      &@               @      �?      @               @      �?       @                      �?      @       @      @                       @       @      @       @                      @      �?      @      �?      @               @      �?       @      �?                       @              �?      6@      :@      "@      �?              �?      "@              *@      9@      $@      0@      @      0@      @      &@      @      @              @      @                       @              @      @              @      "@      �?      "@      �?                      "@       @              R@     �v@      .@      ,@      ,@      @      @      @      @      �?       @      �?              �?       @              @                      @       @              �?      @      �?      �?      �?                      �?              @     �L@     �u@      @@     �s@      1@     Pp@      1@     @m@       @      @       @                      @      .@     �l@      $@      ^@             �H@      $@     �Q@      @              @     �Q@              ?@      @      D@      @      1@      @       @      @                       @       @      .@              &@       @      @       @                      @      �?      7@              3@      �?      @      �?                      @      @     �[@      �?     �Q@      �?      0@      �?      @      �?                      @              $@             �K@      @      D@       @               @      D@       @       @              @       @      �?       @                      �?              @@              ;@      .@     �L@       @      @@              ,@       @      2@      �?      @               @      �?       @               @      �?              �?      ,@      �?                      ,@      *@      9@      &@       @      @              @       @      @       @              @      @      �?      @                      �?      �?               @      1@       @      @      �?              �?      @              @      �?                      *@      9@      >@      9@      4@      4@      4@      (@      4@      (@      ,@      �?      @      �?      @              @      �?      �?              �?      �?                      @      &@      @              �?      &@      @              �?      &@      @      @      @               @      @      @      @                      @      @                      @       @              @                      $@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJW:+LhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKh~�BH4         Z                   �`@�#i����?�           ��@                           �?p�L���?�            `s@              
             �?����X�?             <@������������������������       �                     4@������������������������       �                      @       !       
             �?&Eȧ��?�            �q@              	          ����?�ݏ^���?             �F@                           �?z�G�z�?             4@	                           �?�<ݚ�?             2@
                          �]@�q�q�?             @������������������������       �                     @                           a@�q�q�?             @������������������������       �                      @������������������������       �                     �?                          �]@r�q��?             (@������������������������       �                      @                            K@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @                           �? �o_��?             9@                           �?և���X�?
             ,@������������������������       �                     @                          �^@���!pc�?             &@������������������������       �                     @                          p`@���Q��?             @������������������������       �                     @������������������������       �                      @                           �?�C��2(�?	             &@������������������������       �                     @                            �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @"       7                    �?\ ���?�            �m@#       0                    �?L=�m��?'            �N@$       %                   �k@ףp=
�?#             I@������������������������       �                     A@&       -                    �?     ��?             0@'       (                   �_@�����H�?             "@������������������������       �                     @)       ,       	          @33�?      �?             @*       +                    �O@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @.       /                    @L@և���X�?             @������������������������       �                     @������������������������       �                     @1       6                   �q@�eP*L��?             &@2       3                    �?      �?              @������������������������       �                     @4       5                    \@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @8       M       	          ����?P�9�׸?u             f@9       L                    �?�^����?*            �M@:       ;       	          ����?8��8���?"             H@������������������������       �                     "@<       G                   �[@:�&���?            �C@=       >       	          hff�?�q�q�?	             (@������������������������       �                      @?       F                   �Z@�z�G��?             $@@       E                   �`@      �?              @A       D                   l@      �?             @B       C                   �X@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @H       I                    �?�>����?             ;@������������������������       �                     6@J       K                   �`@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     &@N       Y                   �_@�T�~~4�?K            @]@O       X       	          033@�����?             5@P       W       	          ����?P���Q�?             4@Q       R       	          ����?r�q��?             @������������������������       �                     �?S       V                    \@z�G�z�?             @T       U                   �n@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        
             ,@������������������������       �                     �?������������������������       �        ;             X@[       �                    �?������?
           �z@\       �       	          ��� @���!�=�?�            �n@]       �       	          033�?�W�a=�?�            �l@^       m       
             �?�g�A�E�?~            �i@_       l                    �?��˼��?h             e@`       k                   �t@(;L]n�?I             ^@a       f                    @L@P����?H            �]@b       e                   @[@�K}��?=            �Y@c       d                    c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        ;             Y@g       j                    �L@      �?             0@h       i                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �                      @������������������������       �                    �H@n       �                    �?���"͏�?            �B@o       v       	          ����?�n`���?             ?@p       u                   �p@���|���?             &@q       r                    �?z�G�z�?             @������������������������       �                      @s       t                   �m@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @w       �                   �d@ףp=
�?             4@x       y                   �f@�<ݚ�?             "@������������������������       �                     �?z       {       	          ����?      �?              @������������������������       �                     @|       }                    �G@�q�q�?             @������������������������       �                     �?~                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@�       �                    �?      �?             @�       �       	             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    i@�q�q�?             8@�       �       
             �?����X�?             @������������������������       �                     �?�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   hq@@�0�!��?             1@������������������������       �                     (@�       �                    �?���Q��?             @�       �                   `]@�q�q�?             @������������������������       �                     �?�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?      �?
             0@������������������������       �                     &@�       �                    `@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?(����7�?q            @f@�       �       	          ����?X�<ݚ�?Z             b@�       �                   pn@�;_��?G            @\@�       �                   �e@     ��?"             H@�       �       	             �?�	j*D�?             *@�       �                   �\@X�<ݚ�?             "@������������������������       �                     @�       �                   �c@�q�q�?             @�       �                    d@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   @d@b�h�d.�?            �A@�       �                    �D@d}h���?             <@������������������������       �                      @�       �                   �b@8�Z$���?             :@�       �                   �b@�㙢�c�?             7@�       �       	          ����?��S�ۿ?             .@������������������������       �                     &@�       �                    l@      �?             @������������������������       �                     @������������������������       �                     �?�       �       	          ����?      �?              @�       �                   �b@����X�?             @������������������������       �                     �?�       �                    �?r�q��?             @�       �                   d@      �?             @������������������������       �                     �?�       �       	             �?�q�q�?             @�       �                     J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �L@� ���?%            @P@�       �       
             �?\X��t�?             G@�       �                    �I@HP�s��?             9@������������������������       �                     2@�       �       	          @33�?����X�?             @�       �                   �b@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �       	          ����?؇���X�?             5@�       �                    �?��S�ۿ?
             .@������������������������       �                     &@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @�       �       	          ����?�S����?             3@�       �                   �s@�q�q�?             @�       �                   f@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   �u@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?�       �                   �d@`Jj��?             ?@�       �                   g@XB���?             =@�       �       
             �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     6@�       �                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          833�?�t����?             A@�       �                   ``@      �?              @�       �       	          ����?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �                   pb@ ��WV�?             :@������������������������       �                     5@�       �                   c@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�t�b��)     h�h(h+K ��h-��R�(KK�KK��h_�B�       `u@     �x@     �O@     �n@      4@       @      4@                       @     �E@     �m@      7@      6@      0@      @      ,@      @      @       @      @              �?       @               @      �?              $@       @       @               @       @       @                       @       @              @      2@      @       @      @              @       @              @      @       @      @                       @      �?      $@              @      �?      @      �?                      @      4@      k@      &@      I@      @     �F@              A@      @      &@      �?       @              @      �?      @      �?      �?              �?      �?                       @      @      @              @      @              @      @      @      @              @      @       @               @      @              @              "@     �d@      @      J@      @     �D@              "@      @      @@      @      @       @              @      @      �?      @      �?      @      �?      �?      �?                      �?               @              @       @               @      9@              6@       @      @       @                      @              &@       @     �\@       @      3@      �?      3@      �?      @              �?      �?      @      �?       @      �?                       @               @              ,@      �?                      X@     pq@      b@     `j@     �A@      j@      5@      h@      *@     �d@      @      ]@      @      ]@       @     @Y@      �?      �?      �?              �?      �?              Y@              .@      �?       @      �?              �?       @              *@                       @     �H@              <@      "@      9@      @      @      @      �?      @               @      �?       @      �?                       @      @              2@       @      @       @              �?      @      �?      @               @      �?      �?              �?      �?              �?      �?              &@              @      @      �?      @              @      �?               @              0@       @       @      @      �?              �?      @              @      �?              ,@      @      (@               @      @       @      �?      �?              �?      �?      �?                      �?               @       @      ,@              &@       @      @              @       @              Q@     �[@      P@      T@      O@     �I@     �@@      .@      @      "@      @      @              @      @       @      �?       @      �?                       @      @                      @      =@      @      6@      @               @      6@      @      3@      @      ,@      �?      &@              @      �?      @                      �?      @      @      @       @              �?      @      �?      @      �?      �?               @      �?      �?      �?      �?                      �?      �?               @                      �?      @              @              =@      B@      :@      4@      7@       @      2@              @       @       @       @       @                       @      @              @      2@      �?      ,@              &@      �?      @              @      �?               @      @       @                      @      @      0@       @      @      �?      @              @      �?              �?              �?      (@              (@      �?               @      =@      �?      <@      �?      @      �?                      @              6@      �?      �?      �?                      �?      @      >@      @      @       @      @              @       @              �?              �?      9@              5@      �?      @      �?                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJF<KdhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKŅ�h~�B+         \       
             �?�#i����?�           ��@                           U@4>���?�             u@������������������������       �                     @       '                    �?����s��?�            �t@                           I@��ɶ�"�?�            �i@       	                    �Q@     ��?             0@                          �d@r�q��?             (@������������������������       �                     $@������������������������       �                      @
                           �?      �?             @������������������������       �                     �?������������������������       �                     @       &                    �?�F�l���?y            �g@                          @[@ >�֕�?W            �a@                          `m@���|���?             &@������������������������       �                     @                           @I@և���X�?             @������������������������       �                     @������������������������       �                     @                          pa@0Ƭ!sĮ?Q             `@                           �?@�z�G�?4             T@                           �?@3����?#             K@                          p@ �q�q�?             8@������������������������       �                     4@                          �_@      �?             @                          Pr@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     >@������������������������       �                     :@        %                   �a@��<D�m�?            �H@!       "                    �N@ܷ��?��?             =@������������������������       �                     9@#       $                   @t@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     4@������������������������       �        "            �I@(       S                    �?     x�?L             `@)       F                   �a@Rg��J��?;            �X@*       9       	          ����?և���X�?.            @S@+       8                   �q@�<ݚ�?            �F@,       5                   �c@�p ��?            �D@-       .                   `X@�#-���?            �A@������������������������       �                     �?/       4                   �_@�IєX�?             A@0       3                   �^@8�Z$���?	             *@1       2                    X@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@������������������������       �                     �?������������������������       �                     5@6       7                    h@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @:       E       	          033�?     ��?             @@;       @                    a@PN��T'�?             ;@<       ?                   `@��S�ۿ?             .@=       >                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@A       B                   �c@      �?             (@������������������������       �                     @C       D       	             �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @G       J                    S@�ՙ/�?             5@H       I                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?K       L                    @K@      �?
             0@������������������������       �                     @M       R                   �a@$�q-�?             *@N       Q                    o@r�q��?             @O       P                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @T       U                    d@�r����?             >@������������������������       �        	             .@V       W                    T@������?             .@������������������������       �                      @X       Y                   `r@8�Z$���?             *@������������������������       �                     $@Z       [                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @]       �                    �?L�~m��?           �x@^       �                   �b@`ˡ��Z�?�            Pt@_       v                    �?��c���?�            pq@`       k                   �`@�Z��L��?,            �Q@a       f                     K@ �q�q�?             H@b       c                    �I@؇���X�?             @������������������������       �                     @d       e                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?g       j                   p`@��Y��]�?            �D@h       i                    `@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                     =@l       u                   b@��+7��?             7@m       n                   @g@���Q��?             $@������������������������       �                     @o       p                    �J@�q�q�?             @������������������������       �                     @q       t                    �?�q�q�?             @r       s       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@w       x                   �g@���%�?�             j@������������������������       �        4             S@y       �                   �a@�t:ɨ�?X            �`@z       �                    �?Pq�����?6            @U@{       |                   `h@$�q-�?              J@������������������������       �                     �?}       �                   0i@�IєX�?            �I@~                          �h@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    @K@`�q�0ܴ?            �G@������������������������       �                     >@�       �                    �?�t����?             1@�       �                    _@�r����?
             .@������������������������       �                     @�       �       	             �?�<ݚ�?             "@�       �                   �`@�q�q�?             @������������������������       �                     �?�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                    �@@�       �                    m@`Ql�R�?"            �G@������������������������       �                     7@�       �                   �m@ �q�q�?             8@������������������������       �                     �?������������������������       �                     7@�       �                   Pc@\X��t�?             G@�       �       	          ����?�8��8��?             (@������������������������       �                     @�       �                   @`@z�G�z�?             @�       �                    @B@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �f@�������?             A@�       �                   �l@r٣����?            �@@�       �                   �g@b�2�tk�?
             2@������������������������       �                     $@�       �                   �c@      �?              @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �r@��S�ۿ?
             .@������������������������       �        	             ,@������������������������       �                     �?������������������������       �                     �?�       �                    �?^|�_��?/            �Q@�       �                   �Z@�<ݚ�?             ;@������������������������       �                     @�       �                   �g@      �?             8@�       �                    �G@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �       	          ����?�X�<ݺ?             2@�       �                    a@r�q��?             @������������������������       �                     @�       �                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        
             (@�       �       	          ����?���|���?             F@�       �                    �?�ՙ/�?             5@�       �                   b@������?
             1@�       �                   @]@8�Z$���?             *@�       �                   �a@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �       	             �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    @P@�LQ�1	�?             7@������������������������       �                     4@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�BP       `u@     �x@      q@     �P@              @      q@     �O@     @h@      *@      &@      @      $@       @      $@                       @      �?      @      �?                      @     �f@       @     �`@       @      @      @      @              @      @              @      @             @_@      @     �S@      �?     �J@      �?      7@      �?      4@              @      �?      �?      �?              �?      �?               @              >@              :@              G@      @      :@      @      9@              �?      @      �?                      @      4@             �I@             �S@      I@      J@      G@      F@     �@@     �A@      $@     �A@      @      @@      @              �?      @@       @      &@       @      &@      �?              �?      &@                      �?      5@              @      @              @      @                      @      "@      7@      @      7@      �?      ,@      �?       @               @      �?                      (@      @      "@              @      @       @      @                       @      @               @      *@      @      �?      @                      �?      @      (@      @              �?      (@      �?      @      �?      �?      �?                      �?              @              @      :@      @      .@              &@      @               @      &@       @      $@              �?       @      �?                       @     �Q@     `t@     �@@     @r@      *@     �p@       @     �O@       @      G@      �?      @              @      �?       @               @      �?              �?      D@      �?      &@              &@      �?                      =@      @      1@      @      @      @               @      @              @       @      �?      �?      �?              �?      �?              �?                      *@      @     `i@              S@      @     �_@      @     @T@      @      H@      �?              @      H@      �?      @              @      �?               @     �F@              >@       @      .@       @      *@              @       @      @       @      �?      �?              �?      �?              �?      �?                      @               @             �@@      �?      G@              7@      �?      7@      �?                      7@      4@      :@      &@      �?      @              @      �?      �?      �?              �?      �?              @              "@      9@       @      9@      @      &@              $@      @      �?       @      �?              �?       @              @              �?      ,@              ,@      �?              �?             �B@      A@      5@      @              @      5@      @      @       @      @                       @      1@      �?      @      �?      @               @      �?              �?       @              (@              0@      <@      *@       @      *@      @      &@       @      @       @      @                       @      @               @       @       @                       @              @      @      4@              4@      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJؽ�hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK�h~�B�4         V                    �?�/�$�y�?�           ��@              
             �?�V��Q�?�            0s@       
                    @L@��.N"Ҭ?|            �i@       	                    �? J���#�?f             f@                          h@�K}��?<            �Y@������������������������       �        :            �X@                           d@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        *            �R@              	          @33�?�חF�P�?             ?@                           �?ܷ��?��?             =@                          Ps@��2(&�?             6@                          �O@�����?             5@                           �?z�G�z�?             @������������������������       �                     @                          `_@      �?              @������������������������       �                     �?������������������������       �                     �?                          �_@      �?             0@                           @M@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@������������������������       �                     �?������������������������       �                     @������������������������       �                      @       I                    �?
�c�Z�?B             Y@       "       	          ����?ڤ���?4            @T@       !                    @M@�IєX�?             1@                            @K@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@#       (                    @E@     ��?,             P@$       '                    �?z�G�z�?             @%       &                    �B@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @)       F                    �Q@0B��D�?'            �M@*       1                    �?4և����?%             L@+       0                   �o@���Q��?	             .@,       /                    h@؇���X�?             @-       .                   `[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @2       ?       	          ����?��r._�?            �D@3       8                    �?ҳ�wY;�?             1@4       5       	          ����?z�G�z�?             @������������������������       �                     @6       7                     K@      �?              @������������������������       �                     �?������������������������       �                     �?9       >                   �d@�q�q�?	             (@:       ;                     L@�z�G��?             $@������������������������       �                     @<       =       	          ����?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @@       A                    �N@ �q�q�?             8@������������������������       �                     2@B       C                   �_@r�q��?             @������������������������       �                     @D       E                   Pn@�q�q�?             @������������������������       �                     �?������������������������       �                      @G       H       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @J       U       	             �?�\��N��?             3@K       P                    n@�θ�?	             *@L       M                    �G@�q�q�?             @������������������������       �                     �?N       O                    g@      �?              @������������������������       �                     �?������������������������       �                     �?Q       T                    �?ףp=
�?             $@R       S                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @W       �                   �c@GI2�J�?           �z@X       i                   f@pH?�U��?�            �v@Y       b       	          ����?�8���?H             ]@Z       ]                   �]@PN��T'�?             ;@[       \       
             �?�z�G��?             $@������������������������       �                     @������������������������       �                     @^       a       
             �?�IєX�?	             1@_       `                    @H@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     (@c       d                    @M@�x�E~�?8            @V@������������������������       �                    �C@e       f                   P`@`2U0*��?              I@������������������������       �                    �C@g       h                   a@"pc�
�?             &@������������������������       �                      @������������������������       �                     "@j       �                    �?�qb���?�            `o@k       �       	          033�?<SvLB�?6             W@l       y                   `@� ���?(            @P@m       n                   �Y@����e��?            �@@������������������������       �                     @o       x                    �?�q�q�?             >@p       w       
             �?\X��t�?             7@q       r                   �n@����X�?	             ,@������������������������       �                      @s       v       	          @33�?�q�q�?             @t       u                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     "@������������������������       �                     @z       �       	          ����?     ��?             @@{       �                   �\@      �?             0@|                          �k@r�q��?             @}       ~       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �F@�z�G��?             $@������������������������       �                     �?�       �                   0l@�<ݚ�?             "@������������������������       �                     @�       �                   @e@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                     P@      �?
             0@������������������������       �                     &@�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�����H�?             ;@�       �                    �?�nkK�?             7@������������������������       �        	             2@�       �       	          `ff@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �       	          ����?      �?             @������������������������       �                     �?�       �       	          ���@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �R@0��_��?i            �c@�       �                    t@`1�=7q�?h            �c@�       �                    �J@D��*�4�?[            @a@�       �                    @J@r�q��?             H@�       �                    �?,���i�?            �D@�       �       
             �?��-�=��?            �C@�       �                    @E@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   pb@�L���?            �B@�       �       	          ����? >�֕�?            �A@�       �                    @H@؇���X�?	             ,@�       �                   `c@      �?              @�       �                   p@�q�q�?             @�       �                    �F@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     5@�       �                    �C@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    ]@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                   �[@����?�?<            �V@�       �       	             �?z�G�z�?             @������������������������       �                      @�       �                   �k@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       	             �?`��>�ϗ?9            @U@�       �                   `^@P���Q�?             4@�       �                     N@�����H�?             "@������������������������       �                     @�       �                    \@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             &@������������������������       �        )            @P@�       �                   �t@�S����?             3@�       �                   `\@���Q��?             @������������������������       �                      @�       �                   �e@�q�q�?             @������������������������       �                     �?�       �       	          @33�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             ,@������������������������       �                      @�       �                    �?      �?*             N@�       �       
             �?���Q��?"             I@�       �                    �L@<ݚ)�?             B@�       �                    �?z�G�z�?             >@�       �                   �b@����X�?             5@�       �       	          033�?      �?             4@�       �                   @d@      �?
             0@�       �                    �J@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @I@@4և���?             ,@������������������������       �                     &@�       �                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     "@�       �                   �a@r�q��?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �d@X�Cc�?
             ,@�       �                   Pp@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   `]@�����H�?             "@�       �       	          @33�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KK�KK��h_�B        t@     �y@     �l@     @S@      i@      @     �e@      �?     @Y@      �?     �X@              @      �?      @                      �?     �R@              :@      @      :@      @      3@      @      3@       @      @      �?      @              �?      �?              �?      �?              .@      �?      @      �?              �?      @              (@                      �?      @                       @      =@     �Q@      4@     �N@      �?      0@      �?      @              @      �?                      "@      3@     �F@      @      �?      �?      �?              �?      �?              @              .@      F@      *@     �E@      @      "@      @      �?      �?      �?              �?      �?              @                       @      @      A@      @      &@      �?      @              @      �?      �?      �?                      �?      @      @      @      @              @      @      @      @                      @       @              �?      7@              2@      �?      @              @      �?       @      �?                       @       @      �?              �?       @              "@      $@      @      $@       @      �?      �?              �?      �?              �?      �?              �?      "@      �?       @      �?                       @              @      @             �V@     u@      N@     0s@      @     �[@      @      7@      @      @      @                      @      �?      0@      �?      @              @      �?                      (@       @     �U@             �C@       @      H@             �C@       @      "@       @                      "@      K@     �h@     �C@     �J@      B@      =@      *@      4@      @              $@      4@      $@      *@      $@      @       @               @      @       @      �?              �?       @                      @              "@              @      7@      "@       @       @      �?      @      �?       @      �?                       @              @      @      @              �?      @       @      @              �?       @               @      �?              .@      �?      &@              @      �?      @                      �?      @      8@      �?      6@              2@      �?      @              @      �?               @       @              �?       @      �?       @                      �?      .@      b@      *@      b@      $@      `@       @      D@      @      B@      @     �A@      �?      �?              �?      �?              @      A@       @     �@@       @      (@       @      @       @      @       @      �?              �?       @                      @               @              @              5@      �?      �?              �?      �?              �?      �?      �?                      �?      @      @      @                      @       @      V@      �?      @               @      �?       @      �?                       @      �?      U@      �?      3@      �?       @              @      �?       @               @      �?                      &@             @P@      @      0@      @       @       @              �?       @              �?      �?      �?      �?                      �?              ,@       @              >@      >@      >@      4@      9@      &@      8@      @      .@      @      .@      @      ,@       @      �?      �?              �?      �?              *@      �?      &@               @      �?       @                      �?      �?      @      �?                      @              �?      "@              �?      @              @      �?       @      �?                       @      @      "@      @      �?      @                      �?      �?       @      �?       @               @      �?                      @              $@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJX��vhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKǅ�h~�B�+         N       
             �?���
%�?�           ��@       ;                    �?�˱��H�?�            �r@              	             ���k�c��?�            `o@������������������������       �                      @       &                    �L@�5U��K�?�             o@       #                   h@�X�<ݺ?            �h@                          @\@ؗp�'ʸ?}            �h@                          �q@H�V�e��?             A@	       
                    �E@ܷ��?��?             =@������������������������       �                     *@                           �G@     ��?             0@                          pb@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     $@                           �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @                          �O@@3����?h            @d@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                          �f@��z*�o�?f            �c@                           _@@�`%���?]            `b@                           @L@ �Jj�G�?            �K@������������������������       �                     K@������������������������       �                     �?������������������������       �        >             W@                           �?�8��8��?	             (@������������������������       �                     @       "                    �?z�G�z�?             @        !                   �f@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @$       %                   pn@      �?              @������������������������       �                     �?������������������������       �                     �?'       0                   �`@d,���O�?%            �I@(       /       	          ����?�q�q�?             8@)       .                    �N@@�0�!��?
             1@*       -                   8q@�q�q�?             "@+       ,       	          ����?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @1       :                   @t@�����H�?             ;@2       3                   �a@$�q-�?             :@������������������������       �                     2@4       5                    X@      �?              @������������������������       �                     �?6       7                   0p@؇���X�?             @������������������������       �                     @8       9                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?<       C                   �j@
j*D>�?             J@=       B       	          033�?H%u��?             9@>       ?                    �M@�8��8��?             8@������������������������       �                     ,@@       A                    @N@z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     �?D       G                   �^@l��
I��?             ;@E       F                    �?$�q-�?             *@������������������������       �                     (@������������������������       �                     �?H       K       	          ����?      �?
             ,@I       J                    �?      �?              @������������������������       �                     @������������������������       �                      @L       M                   �]@r�q��?             @������������������������       �                     �?������������������������       �                     @O       �                   �c@ ��7E��?           �z@P       �                   �`@D�qJ�M�?�             x@Q       ~                    �?�Uu� �?q            �g@R       U                    �?p=
ףp�?`             d@S       T                   �_@      �?             @������������������������       �                     @������������������������       �                     @V       W       	          ����?@4և���?\            @c@������������������������       �                    �C@X       Y       	          833�?t��%�?E            �\@������������������������       �                     �?Z       c                    �?x�}b~|�?D            �\@[       `                    �?R���Q�?
             4@\       _                   `o@���Q��?             @]       ^                    `@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?a       b                   Xq@��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?d       e                   @R@heu+��?:            �W@������������������������       �                     �?f       w                    @O@`Jj��?9            @W@g       t       	          033@xL��N�?-            �R@h       i                   �U@      �?(             P@������������������������       �                     �?j       s                    �? ������?'            �O@k       l                   0a@`Ql�R�?            �G@������������������������       �                     B@m       n                   �l@�C��2(�?             &@������������������������       �                     @o       p                    �?r�q��?             @������������������������       �                     @q       r                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     0@u       v                   0m@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@x       }       	             �?�S����?             3@y       z       	          033�?�q�q�?             "@������������������������       �                     @{       |                   �^@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@       �                    �?����"�?             =@�       �                    @E@@�0�!��?
             1@������������������������       �                      @�       �                    �?��S�ۿ?	             .@������������������������       �                     $@�       �                    b@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   �s@�q�q�?             (@�       �                   h@z�G�z�?             $@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    �R@��I�~R�?�            �h@�       �                   �b@؅&�>��?�            `h@�       �                   pb@�}�+r��?V            �`@�       �                   �b@�]��?D            �Y@�       �                    �?��F�D�?A            �X@�       �                    �?`2U0*��?              I@������������������������       �                     (@�       �                    �?�}�+r��?             C@�       �                   �j@��S�ۿ?             >@������������������������       �        	             .@�       �                    �?�r����?
             .@�       �                    l@�8��8��?             (@������������������������       �                     @�       �                    ]@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �        !            �H@�       �                   �j@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?ףp=
�?             >@�       �                    �?�S����?             3@�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �N@؇���X�?             ,@�       �                   �n@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     &@������������������������       �        *             O@������������������������       �                      @�       �                   `l@k��9�?            �F@�       �                   `Y@���|���?             6@������������������������       �                      @�       �                    �?�z�G��?             4@�       �                   �e@@4և���?	             ,@������������������������       �                     (@�       �                    �I@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �J@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?��<b���?             7@�       �                    �B@�8��8��?	             (@������������������������       �                     �?������������������������       �                     &@�       �                   �e@���|���?             &@�       �                    z@�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK�KK��h_�Bp       0s@     �z@     �n@      L@      l@      :@               @      l@      8@     `g@      &@     @g@      $@      ;@      @      :@      @      *@              *@      @      @      @      @                      @      $@              �?      @      �?                      @     �c@      @       @      �?       @                      �?     �c@       @     @b@      �?      K@      �?      K@                      �?      W@              &@      �?      @              @      �?       @      �?              �?       @               @              �?      �?      �?                      �?      C@      *@      ,@      $@      ,@      @      @      @      @      �?      @                      �?               @       @                      @      8@      @      8@       @      2@              @       @              �?      @      �?      @              �?      �?              �?      �?                      �?      6@      >@      @      6@       @      6@              ,@       @       @       @                       @      �?              3@       @      (@      �?      (@                      �?      @      @       @      @              @       @              @      �?              �?      @              N@     0w@     �D@     �u@      @@     �c@      ,@     @b@      @      @              @      @              &@     �a@             �C@      &@      Z@      �?              $@      Z@      @      1@       @      @      �?      @              @      �?              �?              �?      ,@              ,@      �?              @     �U@      �?              @     �U@      @     �Q@       @      O@      �?              �?      O@      �?      G@              B@      �?      $@              @      �?      @              @      �?      �?      �?                      �?              0@      �?      "@      �?                      "@      @      0@      @      @              @      @      �?              �?      @                      $@      2@      &@      ,@      @               @      ,@      �?      $@              @      �?      @                      �?      @       @       @       @       @       @       @                       @              @       @              "@     �g@      @     �g@      @     �_@      @     �X@       @     @X@       @      H@              (@       @      B@       @      <@              .@       @      *@      �?      &@              @      �?      @      �?                      @      �?       @               @      �?                       @             �H@       @       @               @       @              @      ;@      @      0@      �?      @              @      �?               @      (@       @      @       @                      @               @              &@              O@       @              3@      :@      ,@       @               @      ,@      @      *@      �?      (@              �?      �?      �?                      �?      �?      @              @      �?              @      2@      �?      &@      �?                      &@      @      @      @      @              @      @              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���EhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKŅ�h~�B+         ^       	          033�?�r,��?�           ��@       ;       
             �?H;N	�	�?�             x@                          @E@8Ӈ���?�            `p@                          @^@8�A�0��?             6@������������������������       �                     @                          `V@���Q��?             .@������������������������       �                      @       	                    �J@��
ц��?
             *@������������������������       �                     @
                          �]@      �?              @������������������������       �                     @                          `_@���Q��?             @������������������������       �                      @������������������������       �                     @                           �L@��(\���?�             n@                          �q@���fG��?x             f@                           f@@m����?g            �b@������������������������       �        R            �^@                          0f@$�q-�?             :@������������������������       �                     �?                          @b@`2U0*��?             9@������������������������       �                     8@������������������������       �                     �?                          @g@@4և���?             <@                           �? 7���B�?             ;@������������������������       �                     4@                           ]@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?       *                    �?�<ݚ�?%            �O@        !                    `@�t����?             A@������������������������       �                     *@"       #                   �`@��s����?             5@������������������������       �                     �?$       )                   �t@R���Q�?             4@%       &                   d@�KM�]�?             3@������������������������       �        	             ,@'       (                   Pe@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?+       8                    �?J�8���?             =@,       5                    e@�X����?             6@-       0                    ]@�<ݚ�?             2@.       /                   @Z@      �?             @������������������������       �                     �?������������������������       �                     @1       4       	          ����?@4և���?             ,@2       3                   �c@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                      @6       7                   f@      �?             @������������������������       �                     @������������������������       �                     �?9       :                    �?և���X�?             @������������������������       �                     @������������������������       �                     @<       K       	          ����?�&�5y�?J             _@=       B                    �?�m(�X�?4            @U@>       ?                   �d@�J�T�?)            �Q@������������������������       �        '            �P@@       A                   0e@      �?             @������������������������       �                      @������������������������       �                      @C       J                    �?X�Cc�?             ,@D       I                   �q@X�<ݚ�?             "@E       H                    �?r�q��?             @F       G                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @L       [                    �?�	j*D�?            �C@M       P       	          833�?�'�`d�?            �@@N       O                    @K@���Q��?             $@������������������������       �                     @������������������������       �                     @Q       R                    ]@�LQ�1	�?             7@������������������������       �                     �?S       Z                    �?�C��2(�?             6@T       U                   �l@�KM�]�?
             3@������������������������       �                     &@V       W                   �b@      �?              @������������������������       �                     �?X       Y                   0m@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @\       ]                   @j@r�q��?             @������������������������       �                     @������������������������       �                     �?_       �                   �b@д>��C�?�            �u@`       �                   P`@܍�l�p�?�             r@a       �                    �?�P��G7�?Q            @]@b       c                   �U@�	��)��?I            �Y@������������������������       �                     �?d       �                    �?L紂P�?H            �Y@e       h       
             �?��W��?7            @R@f       g                    �N@�q�q�?             @������������������������       �                      @������������������������       �                     �?i       z                   `_@b�h�d.�?4            �Q@j       w       	          033@      �?#             H@k       v                   �m@�����?             E@l       m                    �?�㙢�c�?             7@������������������������       �                     �?n       u                   �m@��2(&�?             6@o       p                    @L@�����?             5@������������������������       �        
             ,@q       t       	          033@����X�?             @r       s                   �\@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     3@x       y                    �J@�q�q�?             @������������������������       �                      @������������������������       �                     @{       |                   �_@���!pc�?             6@������������������������       �                     @}       �       	          033�?�S����?             3@~                           �?      �?              @������������������������       �                      @�       �                   �Y@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             &@������������������������       �                     =@�       �                   �`@և���X�?             ,@������������������������       �                     @�       �                   n@      �?              @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?Pt�nٔ�?e            �e@�       �                    @N@�g<a�?Z            @c@�       �                   P`@`��F:u�?2            �U@������������������������       �                      O@�       �                     M@�J�4�?             9@�       �                   pv@���N8�?             5@������������������������       �                     4@������������������������       �                     �?�       �       
             �?      �?             @������������������������       �                      @�       �                    �M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        (            �P@�       �                    �?���y4F�?             3@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                     K@      �?	             0@�       �                    �?      �?             @������������������������       �                     �?�       �                    b@�q�q�?             @������������������������       �                     �?�       �                   �p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@�       �                    �L@      �?&             M@�       �                    U@P����?             C@������������������������       �                     @�       �       	          ����?����X�?            �A@�       �                   �c@�z�G��?             $@������������������������       �                     @�       �       
             �?���Q��?             @������������������������       �                     �?�       �                   �d@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?H%u��?             9@�       �                    @B@r�q��?             2@������������������������       �                     �?�       �                    �?�t����?             1@������������������������       �                     $@�       �                    �F@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �P@z�G�z�?             4@�       �                    �?      �?
             0@������������������������       �                     @�       �       	          ����?�����H�?             "@�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   Pa@      �?             @������������������������       �                     �?������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�BP       �t@     Py@     �p@     @]@     `m@      ;@      *@      "@      @              @      "@               @      @      @              @      @       @      @              @       @               @      @             �k@      2@     �e@      @     `b@       @     �^@              8@       @              �?      8@      �?      8@                      �?      :@       @      :@      �?      4@              @      �?              �?      @                      �?     �H@      ,@      >@      @      *@              1@      @              �?      1@      @      1@       @      ,@              @       @               @      @                      �?      3@      $@      .@      @      ,@      @      �?      @      �?                      @      *@      �?      &@      �?      &@                      �?       @              �?      @              @      �?              @      @      @                      @      A@     �V@      @     �S@       @     @Q@             �P@       @       @       @                       @      @      "@      @      @      @      �?       @      �?       @                      �?      @                      @              @      ;@      (@      :@      @      @      @      @                      @      4@      @              �?      4@       @      1@       @      &@              @       @              �?      @      �?              �?      @              @              �?      @              @      �?              N@      r@      ?@     0p@      7@     �W@      .@      V@      �?              ,@      V@      ,@     �M@       @      �?       @                      �?      (@      M@      @      E@      @      C@      @      3@      �?              @      3@       @      3@              ,@       @      @       @       @       @                       @              @      �?                      3@       @      @       @                      @      @      0@      @              @      0@      @      @       @              �?      @      �?                      @              &@              =@       @      @      @               @      @       @      �?       @                      �?              @       @     �d@      @     �b@      @     �T@              O@      @      5@      �?      4@              4@      �?              @      �?       @              �?      �?              �?      �?                     �P@      @      .@       @      �?       @                      �?       @      ,@       @       @      �?              �?       @              �?      �?      �?      �?                      �?              (@      =@      =@      9@      *@              @      9@      $@      @      @              @      @       @              �?      @      �?      @                      �?      6@      @      .@      @              �?      .@       @      $@              @       @      @                       @      @              @      0@      �?      .@              @      �?       @      �?      �?      �?                      �?              @      @      �?              �?      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ:9)bhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B8*         �                    �?T8���?�           ��@       q                    �?�yZ����?           �z@       b       	          033�?���X�K�?�            �v@       9       
             �?����j��?�            �s@                           �?��X��?�             l@                           �?`�?�?i            �d@                          �g@`2U0*��?K            @_@              	            �? ;=֦��?I            �^@	       
                    �?���1��??            �Z@������������������������       �        #             M@                          `a@@�E�x�?            �H@������������������������       �                     D@                           b@�����H�?             "@������������������������       �                     @                          �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?              	          ����?�r����?
             .@                          �p@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     "@                           �D@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                    �D@       4                   �e@^l��[B�?$             M@       )                    @K@j�q����?              I@       (                    @F@(N:!���?            �A@       !                   �[@����X�?	             ,@                            �?�q�q�?             @������������������������       �                      @������������������������       �                     �?"       '                    ]@"pc�
�?             &@#       &                    �?�q�q�?             @$       %                   pb@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     5@*       3                    @N@�q�q�?             .@+       ,                    X@X�<ݚ�?             "@������������������������       �                      @-       .                    @M@և���X�?             @������������������������       �                     @/       0                   �`@      �?             @������������������������       �                      @1       2                    a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @5       6                   Pf@      �?              @������������������������       �                     @7       8                   l@z�G�z�?             @������������������������       �                     @������������������������       �                     �?:       I                   �h@�ހ��?:            �W@;       D                     L@���B���?             :@<       C                    �?�����?             5@=       >                    �?P���Q�?             4@������������������������       �                     1@?       @       	          @33�?�q�q�?             @������������������������       �                     �?A       B                   d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?E       H                    �?���Q��?             @F       G                   0a@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?J       _                    �?      �?)             Q@K       X                   Pq@�q�q�?             H@L       S                   �b@П[;U��?             =@M       P                    �?      �?             4@N       O                   �m@�q�q�?             @������������������������       �                     @������������������������       �                      @Q       R                    �?@4և���?             ,@������������������������       �        
             *@������������������������       �                     �?T       U       	          ����?�����H�?             "@������������������������       �                     @V       W                   �l@�q�q�?             @������������������������       �                      @������������������������       �                     �?Y       Z       	          433�?�S����?
             3@������������������������       �                     (@[       \       	          ����?և���X�?             @������������������������       �                      @]       ^                   �r@z�G�z�?             @������������������������       �                     @������������������������       �                     �?`       a                   �^@ףp=
�?             4@������������������������       �                      @������������������������       �                     2@c       j                    @H@0,Tg��?             E@d       i                    �?�	j*D�?             *@e       h                    �E@X�<ݚ�?             "@f       g                    h@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @k       l                    l@ 	��p�?             =@������������������������       �        
             2@m       p                    ^@"pc�
�?             &@n       o                    @N@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @r       w       
             �?=��T�?1            �Q@s       t                   �O@ҳ�wY;�?             A@������������������������       �                     $@u       v       	          hff @�8��8��?             8@������������������������       �                     6@������������������������       �                      @x       �       	          `ff@4?,R��?             B@y       z                   �j@l��\��?             A@������������������������       �                     :@{       |                   pm@      �?              @������������������������       �                      @}       �                    �?r�q��?             @~                          8w@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?�s�ۺ�?�             s@�       �                    �R@���:�?�            pp@�       �                   �Z@��E���?�            `p@�       �                   0a@      �?              @������������������������       �                     @������������������������       �                     @�       �       	          ����?������?�            �o@�       �       
             �?�+e�X�?              I@�       �                   @`@�	j*D�?	             *@������������������������       �                      @�       �                    Y@"pc�
�?             &@������������������������       �                     �?�       �                    h@ףp=
�?             $@�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �_@�L���?            �B@������������������������       �                     .@�       �       	          ����?��2(&�?             6@������������������������       �                     2@�       �                   @_@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �b@Xʃ=��?~            �i@�       �                   P`@`����?z            �h@������������������������       �        ^            �c@�       �                    �?��(\���?             D@�       �                   �W@ �Cc}�?             <@�       �                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �G@`2U0*��?             9@�       �                     E@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     6@������������������������       �                     (@�       �                    �F@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                   �a@�>$�*��?            �D@�       �                   @[@������?             >@������������������������       �                      @�       �                    �?d}h���?             <@�       �       
             �?���!pc�?	             6@������������������������       �                     @�       �                   �\@      �?             0@������������������������       �                     �?�       �       	             �?�q�q�?             .@������������������������       �                     @�       �                   �a@r�q��?             (@������������������������       �                      @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    @O@�C��2(�?	             &@������������������������       �                     @�       �                   `b@      �?             @������������������������       �                     @������������������������       �                     �?�t�b��H      h�h(h+K ��h-��R�(KK�KK��h_�B       �t@     @y@     �q@     `b@      p@      Z@     �n@     @R@     �i@      2@      d@      @      ^@      @     �]@      @     �Z@      �?      M@              H@      �?      D@               @      �?      @               @      �?       @                      �?      *@       @      @       @               @      @              "@              �?       @      �?                       @     �D@             �F@      *@     �D@      "@      ?@      @      $@      @      �?       @               @      �?              "@       @      @       @       @       @       @                       @       @              @              5@              $@      @      @      @               @      @      @      @              �?      @               @      �?      �?              �?      �?              @              @      @      @              �?      @              @      �?             �C@     �K@      @      5@       @      3@      �?      3@              1@      �?       @              �?      �?      �?      �?                      �?      �?              @       @      @      �?              �?      @                      �?      A@      A@      0@      @@      *@      0@      @      .@      @       @      @                       @      �?      *@              *@      �?               @      �?      @               @      �?       @                      �?      @      0@              (@      @      @       @              �?      @              @      �?              2@       @               @      2@              &@      ?@      "@      @      @      @      @      �?              �?      @                      @      @               @      ;@              2@       @      "@       @      �?              �?       @                       @      ;@     �E@      6@      (@              $@      6@       @      6@                       @      @      ?@      @      ?@              :@      @      @       @              �?      @      �?       @               @      �?                      @       @             �G@     p@      8@     �m@      7@     �m@      @      @              @      @              3@     `m@      (@      C@      "@      @               @      "@       @              �?      "@      �?      �?      �?      �?                      �?       @              @      A@              .@      @      3@              2@      @      �?      @                      �?      @     �h@      @     @h@             �c@      @     �B@      @      9@       @      �?       @                      �?      �?      8@      �?       @               @      �?                      6@              (@      @      @      @                      @      �?              7@      2@      6@       @               @      6@      @      0@      @      @              $@      @              �?      $@      @              @      $@       @       @               @       @       @                       @      @              �?      $@              @      �?      @              @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�BHzhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKӅ�h~�B(.         b       	          ����?�[��N�?�           ��@       C       
             �?��)��?�            �v@                          `^@0�|#�p�?�            �o@                           �?V������?            �B@       
                    �?���}<S�?             7@                           �?�����H�?             2@������������������������       �                      @       	                   �]@z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     @                           \@X�Cc�?             ,@������������������������       �                     @                          pb@"pc�
�?             &@                          �_@ףp=
�?             $@������������������������       �                     @                           �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?                           �A@��g�?~            @k@                           �?R���Q�?             4@                          �c@�X�<ݺ?
             2@                           �?؇���X�?             @                          Pc@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@������������������������       �                      @       "                    I@�FVQ&�?s            �h@        !       	          ���ٿ���Q��?             @������������������������       �                      @������������������������       �                     @#       B                   �g@�-j'�?p             h@$       1                    �?�F�l���?o            �g@%       ,                    �O@@P���x�?P            �a@&       +                   0c@`��(�?L            �`@'       *                    �G@ 7���B�?!             K@(       )                   �b@؇���X�?	             ,@������������������������       �                     (@������������������������       �                      @������������������������       �                     D@������������������������       �        +            @T@-       0                    �?z�G�z�?             @.       /       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @2       A                    @M@`�H�/��?            �I@3       @                   Pe@4?,R��?             B@4       7                    �D@�FVQ&�?            �@@5       6                   �h@�q�q�?             @������������������������       �                     �?������������������������       �                      @8       ?                    `@(;L]n�?             >@9       :                   �o@�8��8��?             (@������������������������       �                     "@;       >                    �?�q�q�?             @<       =                    _@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     2@������������������������       �                     @������������������������       �                     .@������������������������       �                      @D       K                    �?��>4��?H             \@E       J                   @_@      �?              @F       G                    �F@      �?             @������������������������       �                      @H       I                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @L       S       	          ����?���c���?B             Z@M       N                    `P@�e���@�?2            @S@������������������������       �        -            �Q@O       R                    �?r�q��?             @P       Q                   `a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @T       ]       	          ����?|��?���?             ;@U       V                   �i@�ՙ/�?             5@������������������������       �                     @W       X                    `@և���X�?             ,@������������������������       �                     @Y       Z                    �?z�G�z�?             $@������������������������       �                     @[       \       	          hff�?�q�q�?             @������������������������       �                      @������������������������       �                     �?^       _                   �l@r�q��?             @������������������������       �                     @`       a                     K@      �?              @������������������������       �                     �?������������������������       �                     �?c       �       
             �?ByL5���?�            �v@d       k                   �_@h�����?%             L@e       f                    �?$�q-�?	             *@������������������������       �                     @g       h                   �f@ףp=
�?             $@������������������������       �                     @i       j       	          033�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?l              	          033@�^�����?            �E@m       n                   �\@���� �?            �D@������������������������       �                     @o       x                   @j@���y4F�?             C@p       w                    b@��
ц��?             *@q       v                   0i@�q�q�?             "@r       s       	             �?      �?             @������������������������       �                      @t       u                   �^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @y       ~                   �d@HP�s��?             9@z       {                    �? �q�q�?             8@������������������������       �                     4@|       }                   �r@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �x@ ��om��?�            ps@�       �                    �?ܴD��?�            �r@�       �                   �n@     ��?'             P@�       �                    n@nM`����?             G@�       �                    �?��i#[�?             E@�       �                   �g@D�n�3�?             3@�       �                   @]@      �?              @������������������������       �                     �?�       �       	          `ff@؇���X�?             @������������������������       �                     @�       �                   @L@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �\@"pc�
�?             &@������������������������       �                     �?�       �       	          `ff@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?�       �                   �e@���}<S�?             7@�       �                    �?���7�?             6@������������������������       �                     5@������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    ]@�X�<ݺ?
             2@������������������������       �                     �?������������������������       �        	             1@�       �                    �?4�ԗj�?�            �m@�       �       	          pff�?l�b�G��?n            `e@�       �       	          033�?���(\��?4             T@�       �                   �s@$�q-�?#             J@�       �                    �?��<D�m�?             �H@������������������������       �                     <@�       �                    @G@؇���X�?             5@�       �                    ^@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   Xr@�����H�?             2@�       �                    �L@      �?             0@�       �                   �Z@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�q�q�?             @�       �                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �?�>4և��?             <@�       �                   �^@������?             1@������������������������       �                     $@�       �                    ]@և���X�?             @������������������������       �                     @�       �                   �g@      �?             @������������������������       �                     �?������������������������       �                     @�       �       	          ����?�C��2(�?             &@�       �                   �\@؇���X�?             @�       �                   @\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    _@x��B�R�?:            �V@�       �                    �J@�C��2(�?             6@�       �                     I@z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     (@�       �                    `P@@	tbA@�?-            @Q@������������������������       �        )             P@�       �                    b@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        ,             Q@�       �                   0c@      �?              @�       �                    X@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B0       �s@     Pz@      o@     �]@     �l@      :@      :@      &@      5@       @      0@       @       @               @       @       @                       @      @              @      "@      @               @      "@      �?      "@              @      �?      @      �?                      @      �?             `i@      .@      1@      @      1@      �?      @      �?       @      �?       @                      �?      @              &@                       @     @g@      (@      @       @               @      @             �f@      $@     �f@       @      a@      @     �`@       @      J@       @      (@       @      (@                       @      D@             @T@              @      �?      �?      �?              �?      �?              @              G@      @      ?@      @      ?@       @       @      �?              �?       @              =@      �?      &@      �?      "@               @      �?      �?      �?      �?                      �?      �?              2@                      @      .@                       @      3@     @W@      @      @      �?      @               @      �?      �?      �?                      �?      @              ,@     �V@      �?      S@             �Q@      �?      @      �?       @               @      �?                      @      *@      ,@       @      *@              @       @      @              @       @       @      @              �?       @               @      �?              @      �?      @              �?      �?              �?      �?             @P@     �r@      ?@      9@      �?      (@              @      �?      "@              @      �?      @              @      �?              >@      *@      >@      &@              @      >@       @      @      @      @      @      @      �?       @              �?      �?      �?                      �?              @      @              7@       @      7@      �?      4@              @      �?      @                      �?              �?               @      A@     Pq@      >@     q@      2@      G@      1@      =@      *@      =@      &@       @       @      @      �?              �?      @              @      �?       @      �?                       @      "@       @              �?      "@      �?      "@                      �?       @      5@      �?      5@              5@      �?              �?              @              �?      1@      �?                      1@      (@     `l@      (@     �c@      "@     �Q@      @      H@      @      G@              <@      @      2@      �?       @      �?                       @       @      0@      �?      .@      �?      @      �?                      @              "@      �?      �?      �?                      �?      �?       @      �?      �?      �?                      �?              �?      @      7@      @      *@              $@      @      @      @              �?      @      �?                      @      �?      $@      �?      @      �?      �?              �?      �?                      @              @      @      V@       @      4@       @       @               @       @                      (@      �?      Q@              P@      �?      @              @      �?                      Q@      @      @      �?      @      �?                      @      @        �t�bubhhubehhub.